magic
tech sky130A
magscale 1 2
timestamp 1640969486
<< error_p >>
rect -653 581 -595 587
rect -461 581 -403 587
rect -269 581 -211 587
rect -77 581 -19 587
rect 115 581 173 587
rect 307 581 365 587
rect 499 581 557 587
rect 691 581 749 587
rect -653 547 -641 581
rect -461 547 -449 581
rect -269 547 -257 581
rect -77 547 -65 581
rect 115 547 127 581
rect 307 547 319 581
rect 499 547 511 581
rect 691 547 703 581
rect -653 541 -595 547
rect -461 541 -403 547
rect -269 541 -211 547
rect -77 541 -19 547
rect 115 541 173 547
rect 307 541 365 547
rect 499 541 557 547
rect 691 541 749 547
rect -749 -547 -691 -541
rect -557 -547 -499 -541
rect -365 -547 -307 -541
rect -173 -547 -115 -541
rect 19 -547 77 -541
rect 211 -547 269 -541
rect 403 -547 461 -541
rect 595 -547 653 -541
rect -749 -581 -737 -547
rect -557 -581 -545 -547
rect -365 -581 -353 -547
rect -173 -581 -161 -547
rect 19 -581 31 -547
rect 211 -581 223 -547
rect 403 -581 415 -547
rect 595 -581 607 -547
rect -749 -587 -691 -581
rect -557 -587 -499 -581
rect -365 -587 -307 -581
rect -173 -587 -115 -581
rect 19 -587 77 -581
rect 211 -587 269 -581
rect 403 -587 461 -581
rect 595 -587 653 -581
<< nwell >>
rect -935 -719 935 719
<< pmos >>
rect -735 -500 -705 500
rect -639 -500 -609 500
rect -543 -500 -513 500
rect -447 -500 -417 500
rect -351 -500 -321 500
rect -255 -500 -225 500
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
rect 225 -500 255 500
rect 321 -500 351 500
rect 417 -500 447 500
rect 513 -500 543 500
rect 609 -500 639 500
rect 705 -500 735 500
<< pdiff >>
rect -797 459 -735 500
rect -797 425 -785 459
rect -751 425 -735 459
rect -797 391 -735 425
rect -797 357 -785 391
rect -751 357 -735 391
rect -797 323 -735 357
rect -797 289 -785 323
rect -751 289 -735 323
rect -797 255 -735 289
rect -797 221 -785 255
rect -751 221 -735 255
rect -797 187 -735 221
rect -797 153 -785 187
rect -751 153 -735 187
rect -797 119 -735 153
rect -797 85 -785 119
rect -751 85 -735 119
rect -797 51 -735 85
rect -797 17 -785 51
rect -751 17 -735 51
rect -797 -17 -735 17
rect -797 -51 -785 -17
rect -751 -51 -735 -17
rect -797 -85 -735 -51
rect -797 -119 -785 -85
rect -751 -119 -735 -85
rect -797 -153 -735 -119
rect -797 -187 -785 -153
rect -751 -187 -735 -153
rect -797 -221 -735 -187
rect -797 -255 -785 -221
rect -751 -255 -735 -221
rect -797 -289 -735 -255
rect -797 -323 -785 -289
rect -751 -323 -735 -289
rect -797 -357 -735 -323
rect -797 -391 -785 -357
rect -751 -391 -735 -357
rect -797 -425 -735 -391
rect -797 -459 -785 -425
rect -751 -459 -735 -425
rect -797 -500 -735 -459
rect -705 459 -639 500
rect -705 425 -689 459
rect -655 425 -639 459
rect -705 391 -639 425
rect -705 357 -689 391
rect -655 357 -639 391
rect -705 323 -639 357
rect -705 289 -689 323
rect -655 289 -639 323
rect -705 255 -639 289
rect -705 221 -689 255
rect -655 221 -639 255
rect -705 187 -639 221
rect -705 153 -689 187
rect -655 153 -639 187
rect -705 119 -639 153
rect -705 85 -689 119
rect -655 85 -639 119
rect -705 51 -639 85
rect -705 17 -689 51
rect -655 17 -639 51
rect -705 -17 -639 17
rect -705 -51 -689 -17
rect -655 -51 -639 -17
rect -705 -85 -639 -51
rect -705 -119 -689 -85
rect -655 -119 -639 -85
rect -705 -153 -639 -119
rect -705 -187 -689 -153
rect -655 -187 -639 -153
rect -705 -221 -639 -187
rect -705 -255 -689 -221
rect -655 -255 -639 -221
rect -705 -289 -639 -255
rect -705 -323 -689 -289
rect -655 -323 -639 -289
rect -705 -357 -639 -323
rect -705 -391 -689 -357
rect -655 -391 -639 -357
rect -705 -425 -639 -391
rect -705 -459 -689 -425
rect -655 -459 -639 -425
rect -705 -500 -639 -459
rect -609 459 -543 500
rect -609 425 -593 459
rect -559 425 -543 459
rect -609 391 -543 425
rect -609 357 -593 391
rect -559 357 -543 391
rect -609 323 -543 357
rect -609 289 -593 323
rect -559 289 -543 323
rect -609 255 -543 289
rect -609 221 -593 255
rect -559 221 -543 255
rect -609 187 -543 221
rect -609 153 -593 187
rect -559 153 -543 187
rect -609 119 -543 153
rect -609 85 -593 119
rect -559 85 -543 119
rect -609 51 -543 85
rect -609 17 -593 51
rect -559 17 -543 51
rect -609 -17 -543 17
rect -609 -51 -593 -17
rect -559 -51 -543 -17
rect -609 -85 -543 -51
rect -609 -119 -593 -85
rect -559 -119 -543 -85
rect -609 -153 -543 -119
rect -609 -187 -593 -153
rect -559 -187 -543 -153
rect -609 -221 -543 -187
rect -609 -255 -593 -221
rect -559 -255 -543 -221
rect -609 -289 -543 -255
rect -609 -323 -593 -289
rect -559 -323 -543 -289
rect -609 -357 -543 -323
rect -609 -391 -593 -357
rect -559 -391 -543 -357
rect -609 -425 -543 -391
rect -609 -459 -593 -425
rect -559 -459 -543 -425
rect -609 -500 -543 -459
rect -513 459 -447 500
rect -513 425 -497 459
rect -463 425 -447 459
rect -513 391 -447 425
rect -513 357 -497 391
rect -463 357 -447 391
rect -513 323 -447 357
rect -513 289 -497 323
rect -463 289 -447 323
rect -513 255 -447 289
rect -513 221 -497 255
rect -463 221 -447 255
rect -513 187 -447 221
rect -513 153 -497 187
rect -463 153 -447 187
rect -513 119 -447 153
rect -513 85 -497 119
rect -463 85 -447 119
rect -513 51 -447 85
rect -513 17 -497 51
rect -463 17 -447 51
rect -513 -17 -447 17
rect -513 -51 -497 -17
rect -463 -51 -447 -17
rect -513 -85 -447 -51
rect -513 -119 -497 -85
rect -463 -119 -447 -85
rect -513 -153 -447 -119
rect -513 -187 -497 -153
rect -463 -187 -447 -153
rect -513 -221 -447 -187
rect -513 -255 -497 -221
rect -463 -255 -447 -221
rect -513 -289 -447 -255
rect -513 -323 -497 -289
rect -463 -323 -447 -289
rect -513 -357 -447 -323
rect -513 -391 -497 -357
rect -463 -391 -447 -357
rect -513 -425 -447 -391
rect -513 -459 -497 -425
rect -463 -459 -447 -425
rect -513 -500 -447 -459
rect -417 459 -351 500
rect -417 425 -401 459
rect -367 425 -351 459
rect -417 391 -351 425
rect -417 357 -401 391
rect -367 357 -351 391
rect -417 323 -351 357
rect -417 289 -401 323
rect -367 289 -351 323
rect -417 255 -351 289
rect -417 221 -401 255
rect -367 221 -351 255
rect -417 187 -351 221
rect -417 153 -401 187
rect -367 153 -351 187
rect -417 119 -351 153
rect -417 85 -401 119
rect -367 85 -351 119
rect -417 51 -351 85
rect -417 17 -401 51
rect -367 17 -351 51
rect -417 -17 -351 17
rect -417 -51 -401 -17
rect -367 -51 -351 -17
rect -417 -85 -351 -51
rect -417 -119 -401 -85
rect -367 -119 -351 -85
rect -417 -153 -351 -119
rect -417 -187 -401 -153
rect -367 -187 -351 -153
rect -417 -221 -351 -187
rect -417 -255 -401 -221
rect -367 -255 -351 -221
rect -417 -289 -351 -255
rect -417 -323 -401 -289
rect -367 -323 -351 -289
rect -417 -357 -351 -323
rect -417 -391 -401 -357
rect -367 -391 -351 -357
rect -417 -425 -351 -391
rect -417 -459 -401 -425
rect -367 -459 -351 -425
rect -417 -500 -351 -459
rect -321 459 -255 500
rect -321 425 -305 459
rect -271 425 -255 459
rect -321 391 -255 425
rect -321 357 -305 391
rect -271 357 -255 391
rect -321 323 -255 357
rect -321 289 -305 323
rect -271 289 -255 323
rect -321 255 -255 289
rect -321 221 -305 255
rect -271 221 -255 255
rect -321 187 -255 221
rect -321 153 -305 187
rect -271 153 -255 187
rect -321 119 -255 153
rect -321 85 -305 119
rect -271 85 -255 119
rect -321 51 -255 85
rect -321 17 -305 51
rect -271 17 -255 51
rect -321 -17 -255 17
rect -321 -51 -305 -17
rect -271 -51 -255 -17
rect -321 -85 -255 -51
rect -321 -119 -305 -85
rect -271 -119 -255 -85
rect -321 -153 -255 -119
rect -321 -187 -305 -153
rect -271 -187 -255 -153
rect -321 -221 -255 -187
rect -321 -255 -305 -221
rect -271 -255 -255 -221
rect -321 -289 -255 -255
rect -321 -323 -305 -289
rect -271 -323 -255 -289
rect -321 -357 -255 -323
rect -321 -391 -305 -357
rect -271 -391 -255 -357
rect -321 -425 -255 -391
rect -321 -459 -305 -425
rect -271 -459 -255 -425
rect -321 -500 -255 -459
rect -225 459 -159 500
rect -225 425 -209 459
rect -175 425 -159 459
rect -225 391 -159 425
rect -225 357 -209 391
rect -175 357 -159 391
rect -225 323 -159 357
rect -225 289 -209 323
rect -175 289 -159 323
rect -225 255 -159 289
rect -225 221 -209 255
rect -175 221 -159 255
rect -225 187 -159 221
rect -225 153 -209 187
rect -175 153 -159 187
rect -225 119 -159 153
rect -225 85 -209 119
rect -175 85 -159 119
rect -225 51 -159 85
rect -225 17 -209 51
rect -175 17 -159 51
rect -225 -17 -159 17
rect -225 -51 -209 -17
rect -175 -51 -159 -17
rect -225 -85 -159 -51
rect -225 -119 -209 -85
rect -175 -119 -159 -85
rect -225 -153 -159 -119
rect -225 -187 -209 -153
rect -175 -187 -159 -153
rect -225 -221 -159 -187
rect -225 -255 -209 -221
rect -175 -255 -159 -221
rect -225 -289 -159 -255
rect -225 -323 -209 -289
rect -175 -323 -159 -289
rect -225 -357 -159 -323
rect -225 -391 -209 -357
rect -175 -391 -159 -357
rect -225 -425 -159 -391
rect -225 -459 -209 -425
rect -175 -459 -159 -425
rect -225 -500 -159 -459
rect -129 459 -63 500
rect -129 425 -113 459
rect -79 425 -63 459
rect -129 391 -63 425
rect -129 357 -113 391
rect -79 357 -63 391
rect -129 323 -63 357
rect -129 289 -113 323
rect -79 289 -63 323
rect -129 255 -63 289
rect -129 221 -113 255
rect -79 221 -63 255
rect -129 187 -63 221
rect -129 153 -113 187
rect -79 153 -63 187
rect -129 119 -63 153
rect -129 85 -113 119
rect -79 85 -63 119
rect -129 51 -63 85
rect -129 17 -113 51
rect -79 17 -63 51
rect -129 -17 -63 17
rect -129 -51 -113 -17
rect -79 -51 -63 -17
rect -129 -85 -63 -51
rect -129 -119 -113 -85
rect -79 -119 -63 -85
rect -129 -153 -63 -119
rect -129 -187 -113 -153
rect -79 -187 -63 -153
rect -129 -221 -63 -187
rect -129 -255 -113 -221
rect -79 -255 -63 -221
rect -129 -289 -63 -255
rect -129 -323 -113 -289
rect -79 -323 -63 -289
rect -129 -357 -63 -323
rect -129 -391 -113 -357
rect -79 -391 -63 -357
rect -129 -425 -63 -391
rect -129 -459 -113 -425
rect -79 -459 -63 -425
rect -129 -500 -63 -459
rect -33 459 33 500
rect -33 425 -17 459
rect 17 425 33 459
rect -33 391 33 425
rect -33 357 -17 391
rect 17 357 33 391
rect -33 323 33 357
rect -33 289 -17 323
rect 17 289 33 323
rect -33 255 33 289
rect -33 221 -17 255
rect 17 221 33 255
rect -33 187 33 221
rect -33 153 -17 187
rect 17 153 33 187
rect -33 119 33 153
rect -33 85 -17 119
rect 17 85 33 119
rect -33 51 33 85
rect -33 17 -17 51
rect 17 17 33 51
rect -33 -17 33 17
rect -33 -51 -17 -17
rect 17 -51 33 -17
rect -33 -85 33 -51
rect -33 -119 -17 -85
rect 17 -119 33 -85
rect -33 -153 33 -119
rect -33 -187 -17 -153
rect 17 -187 33 -153
rect -33 -221 33 -187
rect -33 -255 -17 -221
rect 17 -255 33 -221
rect -33 -289 33 -255
rect -33 -323 -17 -289
rect 17 -323 33 -289
rect -33 -357 33 -323
rect -33 -391 -17 -357
rect 17 -391 33 -357
rect -33 -425 33 -391
rect -33 -459 -17 -425
rect 17 -459 33 -425
rect -33 -500 33 -459
rect 63 459 129 500
rect 63 425 79 459
rect 113 425 129 459
rect 63 391 129 425
rect 63 357 79 391
rect 113 357 129 391
rect 63 323 129 357
rect 63 289 79 323
rect 113 289 129 323
rect 63 255 129 289
rect 63 221 79 255
rect 113 221 129 255
rect 63 187 129 221
rect 63 153 79 187
rect 113 153 129 187
rect 63 119 129 153
rect 63 85 79 119
rect 113 85 129 119
rect 63 51 129 85
rect 63 17 79 51
rect 113 17 129 51
rect 63 -17 129 17
rect 63 -51 79 -17
rect 113 -51 129 -17
rect 63 -85 129 -51
rect 63 -119 79 -85
rect 113 -119 129 -85
rect 63 -153 129 -119
rect 63 -187 79 -153
rect 113 -187 129 -153
rect 63 -221 129 -187
rect 63 -255 79 -221
rect 113 -255 129 -221
rect 63 -289 129 -255
rect 63 -323 79 -289
rect 113 -323 129 -289
rect 63 -357 129 -323
rect 63 -391 79 -357
rect 113 -391 129 -357
rect 63 -425 129 -391
rect 63 -459 79 -425
rect 113 -459 129 -425
rect 63 -500 129 -459
rect 159 459 225 500
rect 159 425 175 459
rect 209 425 225 459
rect 159 391 225 425
rect 159 357 175 391
rect 209 357 225 391
rect 159 323 225 357
rect 159 289 175 323
rect 209 289 225 323
rect 159 255 225 289
rect 159 221 175 255
rect 209 221 225 255
rect 159 187 225 221
rect 159 153 175 187
rect 209 153 225 187
rect 159 119 225 153
rect 159 85 175 119
rect 209 85 225 119
rect 159 51 225 85
rect 159 17 175 51
rect 209 17 225 51
rect 159 -17 225 17
rect 159 -51 175 -17
rect 209 -51 225 -17
rect 159 -85 225 -51
rect 159 -119 175 -85
rect 209 -119 225 -85
rect 159 -153 225 -119
rect 159 -187 175 -153
rect 209 -187 225 -153
rect 159 -221 225 -187
rect 159 -255 175 -221
rect 209 -255 225 -221
rect 159 -289 225 -255
rect 159 -323 175 -289
rect 209 -323 225 -289
rect 159 -357 225 -323
rect 159 -391 175 -357
rect 209 -391 225 -357
rect 159 -425 225 -391
rect 159 -459 175 -425
rect 209 -459 225 -425
rect 159 -500 225 -459
rect 255 459 321 500
rect 255 425 271 459
rect 305 425 321 459
rect 255 391 321 425
rect 255 357 271 391
rect 305 357 321 391
rect 255 323 321 357
rect 255 289 271 323
rect 305 289 321 323
rect 255 255 321 289
rect 255 221 271 255
rect 305 221 321 255
rect 255 187 321 221
rect 255 153 271 187
rect 305 153 321 187
rect 255 119 321 153
rect 255 85 271 119
rect 305 85 321 119
rect 255 51 321 85
rect 255 17 271 51
rect 305 17 321 51
rect 255 -17 321 17
rect 255 -51 271 -17
rect 305 -51 321 -17
rect 255 -85 321 -51
rect 255 -119 271 -85
rect 305 -119 321 -85
rect 255 -153 321 -119
rect 255 -187 271 -153
rect 305 -187 321 -153
rect 255 -221 321 -187
rect 255 -255 271 -221
rect 305 -255 321 -221
rect 255 -289 321 -255
rect 255 -323 271 -289
rect 305 -323 321 -289
rect 255 -357 321 -323
rect 255 -391 271 -357
rect 305 -391 321 -357
rect 255 -425 321 -391
rect 255 -459 271 -425
rect 305 -459 321 -425
rect 255 -500 321 -459
rect 351 459 417 500
rect 351 425 367 459
rect 401 425 417 459
rect 351 391 417 425
rect 351 357 367 391
rect 401 357 417 391
rect 351 323 417 357
rect 351 289 367 323
rect 401 289 417 323
rect 351 255 417 289
rect 351 221 367 255
rect 401 221 417 255
rect 351 187 417 221
rect 351 153 367 187
rect 401 153 417 187
rect 351 119 417 153
rect 351 85 367 119
rect 401 85 417 119
rect 351 51 417 85
rect 351 17 367 51
rect 401 17 417 51
rect 351 -17 417 17
rect 351 -51 367 -17
rect 401 -51 417 -17
rect 351 -85 417 -51
rect 351 -119 367 -85
rect 401 -119 417 -85
rect 351 -153 417 -119
rect 351 -187 367 -153
rect 401 -187 417 -153
rect 351 -221 417 -187
rect 351 -255 367 -221
rect 401 -255 417 -221
rect 351 -289 417 -255
rect 351 -323 367 -289
rect 401 -323 417 -289
rect 351 -357 417 -323
rect 351 -391 367 -357
rect 401 -391 417 -357
rect 351 -425 417 -391
rect 351 -459 367 -425
rect 401 -459 417 -425
rect 351 -500 417 -459
rect 447 459 513 500
rect 447 425 463 459
rect 497 425 513 459
rect 447 391 513 425
rect 447 357 463 391
rect 497 357 513 391
rect 447 323 513 357
rect 447 289 463 323
rect 497 289 513 323
rect 447 255 513 289
rect 447 221 463 255
rect 497 221 513 255
rect 447 187 513 221
rect 447 153 463 187
rect 497 153 513 187
rect 447 119 513 153
rect 447 85 463 119
rect 497 85 513 119
rect 447 51 513 85
rect 447 17 463 51
rect 497 17 513 51
rect 447 -17 513 17
rect 447 -51 463 -17
rect 497 -51 513 -17
rect 447 -85 513 -51
rect 447 -119 463 -85
rect 497 -119 513 -85
rect 447 -153 513 -119
rect 447 -187 463 -153
rect 497 -187 513 -153
rect 447 -221 513 -187
rect 447 -255 463 -221
rect 497 -255 513 -221
rect 447 -289 513 -255
rect 447 -323 463 -289
rect 497 -323 513 -289
rect 447 -357 513 -323
rect 447 -391 463 -357
rect 497 -391 513 -357
rect 447 -425 513 -391
rect 447 -459 463 -425
rect 497 -459 513 -425
rect 447 -500 513 -459
rect 543 459 609 500
rect 543 425 559 459
rect 593 425 609 459
rect 543 391 609 425
rect 543 357 559 391
rect 593 357 609 391
rect 543 323 609 357
rect 543 289 559 323
rect 593 289 609 323
rect 543 255 609 289
rect 543 221 559 255
rect 593 221 609 255
rect 543 187 609 221
rect 543 153 559 187
rect 593 153 609 187
rect 543 119 609 153
rect 543 85 559 119
rect 593 85 609 119
rect 543 51 609 85
rect 543 17 559 51
rect 593 17 609 51
rect 543 -17 609 17
rect 543 -51 559 -17
rect 593 -51 609 -17
rect 543 -85 609 -51
rect 543 -119 559 -85
rect 593 -119 609 -85
rect 543 -153 609 -119
rect 543 -187 559 -153
rect 593 -187 609 -153
rect 543 -221 609 -187
rect 543 -255 559 -221
rect 593 -255 609 -221
rect 543 -289 609 -255
rect 543 -323 559 -289
rect 593 -323 609 -289
rect 543 -357 609 -323
rect 543 -391 559 -357
rect 593 -391 609 -357
rect 543 -425 609 -391
rect 543 -459 559 -425
rect 593 -459 609 -425
rect 543 -500 609 -459
rect 639 459 705 500
rect 639 425 655 459
rect 689 425 705 459
rect 639 391 705 425
rect 639 357 655 391
rect 689 357 705 391
rect 639 323 705 357
rect 639 289 655 323
rect 689 289 705 323
rect 639 255 705 289
rect 639 221 655 255
rect 689 221 705 255
rect 639 187 705 221
rect 639 153 655 187
rect 689 153 705 187
rect 639 119 705 153
rect 639 85 655 119
rect 689 85 705 119
rect 639 51 705 85
rect 639 17 655 51
rect 689 17 705 51
rect 639 -17 705 17
rect 639 -51 655 -17
rect 689 -51 705 -17
rect 639 -85 705 -51
rect 639 -119 655 -85
rect 689 -119 705 -85
rect 639 -153 705 -119
rect 639 -187 655 -153
rect 689 -187 705 -153
rect 639 -221 705 -187
rect 639 -255 655 -221
rect 689 -255 705 -221
rect 639 -289 705 -255
rect 639 -323 655 -289
rect 689 -323 705 -289
rect 639 -357 705 -323
rect 639 -391 655 -357
rect 689 -391 705 -357
rect 639 -425 705 -391
rect 639 -459 655 -425
rect 689 -459 705 -425
rect 639 -500 705 -459
rect 735 459 797 500
rect 735 425 751 459
rect 785 425 797 459
rect 735 391 797 425
rect 735 357 751 391
rect 785 357 797 391
rect 735 323 797 357
rect 735 289 751 323
rect 785 289 797 323
rect 735 255 797 289
rect 735 221 751 255
rect 785 221 797 255
rect 735 187 797 221
rect 735 153 751 187
rect 785 153 797 187
rect 735 119 797 153
rect 735 85 751 119
rect 785 85 797 119
rect 735 51 797 85
rect 735 17 751 51
rect 785 17 797 51
rect 735 -17 797 17
rect 735 -51 751 -17
rect 785 -51 797 -17
rect 735 -85 797 -51
rect 735 -119 751 -85
rect 785 -119 797 -85
rect 735 -153 797 -119
rect 735 -187 751 -153
rect 785 -187 797 -153
rect 735 -221 797 -187
rect 735 -255 751 -221
rect 785 -255 797 -221
rect 735 -289 797 -255
rect 735 -323 751 -289
rect 785 -323 797 -289
rect 735 -357 797 -323
rect 735 -391 751 -357
rect 785 -391 797 -357
rect 735 -425 797 -391
rect 735 -459 751 -425
rect 785 -459 797 -425
rect 735 -500 797 -459
<< pdiffc >>
rect -785 425 -751 459
rect -785 357 -751 391
rect -785 289 -751 323
rect -785 221 -751 255
rect -785 153 -751 187
rect -785 85 -751 119
rect -785 17 -751 51
rect -785 -51 -751 -17
rect -785 -119 -751 -85
rect -785 -187 -751 -153
rect -785 -255 -751 -221
rect -785 -323 -751 -289
rect -785 -391 -751 -357
rect -785 -459 -751 -425
rect -689 425 -655 459
rect -689 357 -655 391
rect -689 289 -655 323
rect -689 221 -655 255
rect -689 153 -655 187
rect -689 85 -655 119
rect -689 17 -655 51
rect -689 -51 -655 -17
rect -689 -119 -655 -85
rect -689 -187 -655 -153
rect -689 -255 -655 -221
rect -689 -323 -655 -289
rect -689 -391 -655 -357
rect -689 -459 -655 -425
rect -593 425 -559 459
rect -593 357 -559 391
rect -593 289 -559 323
rect -593 221 -559 255
rect -593 153 -559 187
rect -593 85 -559 119
rect -593 17 -559 51
rect -593 -51 -559 -17
rect -593 -119 -559 -85
rect -593 -187 -559 -153
rect -593 -255 -559 -221
rect -593 -323 -559 -289
rect -593 -391 -559 -357
rect -593 -459 -559 -425
rect -497 425 -463 459
rect -497 357 -463 391
rect -497 289 -463 323
rect -497 221 -463 255
rect -497 153 -463 187
rect -497 85 -463 119
rect -497 17 -463 51
rect -497 -51 -463 -17
rect -497 -119 -463 -85
rect -497 -187 -463 -153
rect -497 -255 -463 -221
rect -497 -323 -463 -289
rect -497 -391 -463 -357
rect -497 -459 -463 -425
rect -401 425 -367 459
rect -401 357 -367 391
rect -401 289 -367 323
rect -401 221 -367 255
rect -401 153 -367 187
rect -401 85 -367 119
rect -401 17 -367 51
rect -401 -51 -367 -17
rect -401 -119 -367 -85
rect -401 -187 -367 -153
rect -401 -255 -367 -221
rect -401 -323 -367 -289
rect -401 -391 -367 -357
rect -401 -459 -367 -425
rect -305 425 -271 459
rect -305 357 -271 391
rect -305 289 -271 323
rect -305 221 -271 255
rect -305 153 -271 187
rect -305 85 -271 119
rect -305 17 -271 51
rect -305 -51 -271 -17
rect -305 -119 -271 -85
rect -305 -187 -271 -153
rect -305 -255 -271 -221
rect -305 -323 -271 -289
rect -305 -391 -271 -357
rect -305 -459 -271 -425
rect -209 425 -175 459
rect -209 357 -175 391
rect -209 289 -175 323
rect -209 221 -175 255
rect -209 153 -175 187
rect -209 85 -175 119
rect -209 17 -175 51
rect -209 -51 -175 -17
rect -209 -119 -175 -85
rect -209 -187 -175 -153
rect -209 -255 -175 -221
rect -209 -323 -175 -289
rect -209 -391 -175 -357
rect -209 -459 -175 -425
rect -113 425 -79 459
rect -113 357 -79 391
rect -113 289 -79 323
rect -113 221 -79 255
rect -113 153 -79 187
rect -113 85 -79 119
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -119 -79 -85
rect -113 -187 -79 -153
rect -113 -255 -79 -221
rect -113 -323 -79 -289
rect -113 -391 -79 -357
rect -113 -459 -79 -425
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect 79 425 113 459
rect 79 357 113 391
rect 79 289 113 323
rect 79 221 113 255
rect 79 153 113 187
rect 79 85 113 119
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -119 113 -85
rect 79 -187 113 -153
rect 79 -255 113 -221
rect 79 -323 113 -289
rect 79 -391 113 -357
rect 79 -459 113 -425
rect 175 425 209 459
rect 175 357 209 391
rect 175 289 209 323
rect 175 221 209 255
rect 175 153 209 187
rect 175 85 209 119
rect 175 17 209 51
rect 175 -51 209 -17
rect 175 -119 209 -85
rect 175 -187 209 -153
rect 175 -255 209 -221
rect 175 -323 209 -289
rect 175 -391 209 -357
rect 175 -459 209 -425
rect 271 425 305 459
rect 271 357 305 391
rect 271 289 305 323
rect 271 221 305 255
rect 271 153 305 187
rect 271 85 305 119
rect 271 17 305 51
rect 271 -51 305 -17
rect 271 -119 305 -85
rect 271 -187 305 -153
rect 271 -255 305 -221
rect 271 -323 305 -289
rect 271 -391 305 -357
rect 271 -459 305 -425
rect 367 425 401 459
rect 367 357 401 391
rect 367 289 401 323
rect 367 221 401 255
rect 367 153 401 187
rect 367 85 401 119
rect 367 17 401 51
rect 367 -51 401 -17
rect 367 -119 401 -85
rect 367 -187 401 -153
rect 367 -255 401 -221
rect 367 -323 401 -289
rect 367 -391 401 -357
rect 367 -459 401 -425
rect 463 425 497 459
rect 463 357 497 391
rect 463 289 497 323
rect 463 221 497 255
rect 463 153 497 187
rect 463 85 497 119
rect 463 17 497 51
rect 463 -51 497 -17
rect 463 -119 497 -85
rect 463 -187 497 -153
rect 463 -255 497 -221
rect 463 -323 497 -289
rect 463 -391 497 -357
rect 463 -459 497 -425
rect 559 425 593 459
rect 559 357 593 391
rect 559 289 593 323
rect 559 221 593 255
rect 559 153 593 187
rect 559 85 593 119
rect 559 17 593 51
rect 559 -51 593 -17
rect 559 -119 593 -85
rect 559 -187 593 -153
rect 559 -255 593 -221
rect 559 -323 593 -289
rect 559 -391 593 -357
rect 559 -459 593 -425
rect 655 425 689 459
rect 655 357 689 391
rect 655 289 689 323
rect 655 221 689 255
rect 655 153 689 187
rect 655 85 689 119
rect 655 17 689 51
rect 655 -51 689 -17
rect 655 -119 689 -85
rect 655 -187 689 -153
rect 655 -255 689 -221
rect 655 -323 689 -289
rect 655 -391 689 -357
rect 655 -459 689 -425
rect 751 425 785 459
rect 751 357 785 391
rect 751 289 785 323
rect 751 221 785 255
rect 751 153 785 187
rect 751 85 785 119
rect 751 17 785 51
rect 751 -51 785 -17
rect 751 -119 785 -85
rect 751 -187 785 -153
rect 751 -255 785 -221
rect 751 -323 785 -289
rect 751 -391 785 -357
rect 751 -459 785 -425
<< nsubdiff >>
rect -899 649 -799 683
rect -765 649 -731 683
rect -697 649 -663 683
rect -629 649 -595 683
rect -561 649 -527 683
rect -493 649 -459 683
rect -425 649 -391 683
rect -357 649 -323 683
rect -289 649 -255 683
rect -221 649 -187 683
rect -153 649 -119 683
rect -85 649 -51 683
rect -17 649 17 683
rect 51 649 85 683
rect 119 649 153 683
rect 187 649 221 683
rect 255 649 289 683
rect 323 649 357 683
rect 391 649 425 683
rect 459 649 493 683
rect 527 649 561 683
rect 595 649 629 683
rect 663 649 697 683
rect 731 649 765 683
rect 799 649 899 683
rect -899 561 -865 649
rect 865 561 899 649
rect -899 493 -865 527
rect -899 425 -865 459
rect -899 357 -865 391
rect -899 289 -865 323
rect -899 221 -865 255
rect -899 153 -865 187
rect -899 85 -865 119
rect -899 17 -865 51
rect -899 -51 -865 -17
rect -899 -119 -865 -85
rect -899 -187 -865 -153
rect -899 -255 -865 -221
rect -899 -323 -865 -289
rect -899 -391 -865 -357
rect -899 -459 -865 -425
rect -899 -527 -865 -493
rect 865 493 899 527
rect 865 425 899 459
rect 865 357 899 391
rect 865 289 899 323
rect 865 221 899 255
rect 865 153 899 187
rect 865 85 899 119
rect 865 17 899 51
rect 865 -51 899 -17
rect 865 -119 899 -85
rect 865 -187 899 -153
rect 865 -255 899 -221
rect 865 -323 899 -289
rect 865 -391 899 -357
rect 865 -459 899 -425
rect 865 -527 899 -493
rect -899 -649 -865 -561
rect 865 -649 899 -561
rect -899 -683 -799 -649
rect -765 -683 -731 -649
rect -697 -683 -663 -649
rect -629 -683 -595 -649
rect -561 -683 -527 -649
rect -493 -683 -459 -649
rect -425 -683 -391 -649
rect -357 -683 -323 -649
rect -289 -683 -255 -649
rect -221 -683 -187 -649
rect -153 -683 -119 -649
rect -85 -683 -51 -649
rect -17 -683 17 -649
rect 51 -683 85 -649
rect 119 -683 153 -649
rect 187 -683 221 -649
rect 255 -683 289 -649
rect 323 -683 357 -649
rect 391 -683 425 -649
rect 459 -683 493 -649
rect 527 -683 561 -649
rect 595 -683 629 -649
rect 663 -683 697 -649
rect 731 -683 765 -649
rect 799 -683 899 -649
<< nsubdiffcont >>
rect -799 649 -765 683
rect -731 649 -697 683
rect -663 649 -629 683
rect -595 649 -561 683
rect -527 649 -493 683
rect -459 649 -425 683
rect -391 649 -357 683
rect -323 649 -289 683
rect -255 649 -221 683
rect -187 649 -153 683
rect -119 649 -85 683
rect -51 649 -17 683
rect 17 649 51 683
rect 85 649 119 683
rect 153 649 187 683
rect 221 649 255 683
rect 289 649 323 683
rect 357 649 391 683
rect 425 649 459 683
rect 493 649 527 683
rect 561 649 595 683
rect 629 649 663 683
rect 697 649 731 683
rect 765 649 799 683
rect -899 527 -865 561
rect 865 527 899 561
rect -899 459 -865 493
rect -899 391 -865 425
rect -899 323 -865 357
rect -899 255 -865 289
rect -899 187 -865 221
rect -899 119 -865 153
rect -899 51 -865 85
rect -899 -17 -865 17
rect -899 -85 -865 -51
rect -899 -153 -865 -119
rect -899 -221 -865 -187
rect -899 -289 -865 -255
rect -899 -357 -865 -323
rect -899 -425 -865 -391
rect -899 -493 -865 -459
rect 865 459 899 493
rect 865 391 899 425
rect 865 323 899 357
rect 865 255 899 289
rect 865 187 899 221
rect 865 119 899 153
rect 865 51 899 85
rect 865 -17 899 17
rect 865 -85 899 -51
rect 865 -153 899 -119
rect 865 -221 899 -187
rect 865 -289 899 -255
rect 865 -357 899 -323
rect 865 -425 899 -391
rect 865 -493 899 -459
rect -899 -561 -865 -527
rect 865 -561 899 -527
rect -799 -683 -765 -649
rect -731 -683 -697 -649
rect -663 -683 -629 -649
rect -595 -683 -561 -649
rect -527 -683 -493 -649
rect -459 -683 -425 -649
rect -391 -683 -357 -649
rect -323 -683 -289 -649
rect -255 -683 -221 -649
rect -187 -683 -153 -649
rect -119 -683 -85 -649
rect -51 -683 -17 -649
rect 17 -683 51 -649
rect 85 -683 119 -649
rect 153 -683 187 -649
rect 221 -683 255 -649
rect 289 -683 323 -649
rect 357 -683 391 -649
rect 425 -683 459 -649
rect 493 -683 527 -649
rect 561 -683 595 -649
rect 629 -683 663 -649
rect 697 -683 731 -649
rect 765 -683 799 -649
<< poly >>
rect -657 581 -591 597
rect -657 547 -641 581
rect -607 547 -591 581
rect -657 531 -591 547
rect -465 581 -399 597
rect -465 547 -449 581
rect -415 547 -399 581
rect -465 531 -399 547
rect -273 581 -207 597
rect -273 547 -257 581
rect -223 547 -207 581
rect -273 531 -207 547
rect -81 581 -15 597
rect -81 547 -65 581
rect -31 547 -15 581
rect -81 531 -15 547
rect 111 581 177 597
rect 111 547 127 581
rect 161 547 177 581
rect 111 531 177 547
rect 303 581 369 597
rect 303 547 319 581
rect 353 547 369 581
rect 303 531 369 547
rect 495 581 561 597
rect 495 547 511 581
rect 545 547 561 581
rect 495 531 561 547
rect 687 581 753 597
rect 687 547 703 581
rect 737 547 753 581
rect 687 531 753 547
rect -735 500 -705 526
rect -639 500 -609 531
rect -543 500 -513 526
rect -447 500 -417 531
rect -351 500 -321 526
rect -255 500 -225 531
rect -159 500 -129 526
rect -63 500 -33 531
rect 33 500 63 526
rect 129 500 159 531
rect 225 500 255 526
rect 321 500 351 531
rect 417 500 447 526
rect 513 500 543 531
rect 609 500 639 526
rect 705 500 735 531
rect -735 -531 -705 -500
rect -639 -526 -609 -500
rect -543 -531 -513 -500
rect -447 -526 -417 -500
rect -351 -531 -321 -500
rect -255 -526 -225 -500
rect -159 -531 -129 -500
rect -63 -526 -33 -500
rect 33 -531 63 -500
rect 129 -526 159 -500
rect 225 -531 255 -500
rect 321 -526 351 -500
rect 417 -531 447 -500
rect 513 -526 543 -500
rect 609 -531 639 -500
rect 705 -526 735 -500
rect -753 -547 -687 -531
rect -753 -581 -737 -547
rect -703 -581 -687 -547
rect -753 -597 -687 -581
rect -561 -547 -495 -531
rect -561 -581 -545 -547
rect -511 -581 -495 -547
rect -561 -597 -495 -581
rect -369 -547 -303 -531
rect -369 -581 -353 -547
rect -319 -581 -303 -547
rect -369 -597 -303 -581
rect -177 -547 -111 -531
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect -177 -597 -111 -581
rect 15 -547 81 -531
rect 15 -581 31 -547
rect 65 -581 81 -547
rect 15 -597 81 -581
rect 207 -547 273 -531
rect 207 -581 223 -547
rect 257 -581 273 -547
rect 207 -597 273 -581
rect 399 -547 465 -531
rect 399 -581 415 -547
rect 449 -581 465 -547
rect 399 -597 465 -581
rect 591 -547 657 -531
rect 591 -581 607 -547
rect 641 -581 657 -547
rect 591 -597 657 -581
<< polycont >>
rect -641 547 -607 581
rect -449 547 -415 581
rect -257 547 -223 581
rect -65 547 -31 581
rect 127 547 161 581
rect 319 547 353 581
rect 511 547 545 581
rect 703 547 737 581
rect -737 -581 -703 -547
rect -545 -581 -511 -547
rect -353 -581 -319 -547
rect -161 -581 -127 -547
rect 31 -581 65 -547
rect 223 -581 257 -547
rect 415 -581 449 -547
rect 607 -581 641 -547
<< locali >>
rect -899 649 -799 683
rect -765 649 -731 683
rect -697 649 -663 683
rect -629 649 -595 683
rect -561 649 -527 683
rect -493 649 -459 683
rect -425 649 -391 683
rect -357 649 -323 683
rect -289 649 -255 683
rect -221 649 -187 683
rect -153 649 -119 683
rect -85 649 -51 683
rect -17 649 17 683
rect 51 649 85 683
rect 119 649 153 683
rect 187 649 221 683
rect 255 649 289 683
rect 323 649 357 683
rect 391 649 425 683
rect 459 649 493 683
rect 527 649 561 683
rect 595 649 629 683
rect 663 649 697 683
rect 731 649 765 683
rect 799 649 899 683
rect -899 561 -865 649
rect -657 547 -641 581
rect -607 547 -591 581
rect -465 547 -449 581
rect -415 547 -399 581
rect -273 547 -257 581
rect -223 547 -207 581
rect -81 547 -65 581
rect -31 547 -15 581
rect 111 547 127 581
rect 161 547 177 581
rect 303 547 319 581
rect 353 547 369 581
rect 495 547 511 581
rect 545 547 561 581
rect 687 547 703 581
rect 737 547 753 581
rect 865 561 899 649
rect -899 493 -865 527
rect -899 425 -865 459
rect -899 357 -865 391
rect -899 289 -865 323
rect -899 221 -865 255
rect -899 153 -865 187
rect -899 85 -865 119
rect -899 17 -865 51
rect -899 -51 -865 -17
rect -899 -119 -865 -85
rect -899 -187 -865 -153
rect -899 -255 -865 -221
rect -899 -323 -865 -289
rect -899 -391 -865 -357
rect -899 -459 -865 -425
rect -899 -527 -865 -493
rect -785 485 -751 504
rect -785 413 -751 425
rect -785 341 -751 357
rect -785 269 -751 289
rect -785 197 -751 221
rect -785 125 -751 153
rect -785 53 -751 85
rect -785 -17 -751 17
rect -785 -85 -751 -53
rect -785 -153 -751 -125
rect -785 -221 -751 -197
rect -785 -289 -751 -269
rect -785 -357 -751 -341
rect -785 -425 -751 -413
rect -785 -504 -751 -485
rect -689 485 -655 504
rect -689 413 -655 425
rect -689 341 -655 357
rect -689 269 -655 289
rect -689 197 -655 221
rect -689 125 -655 153
rect -689 53 -655 85
rect -689 -17 -655 17
rect -689 -85 -655 -53
rect -689 -153 -655 -125
rect -689 -221 -655 -197
rect -689 -289 -655 -269
rect -689 -357 -655 -341
rect -689 -425 -655 -413
rect -689 -504 -655 -485
rect -593 485 -559 504
rect -593 413 -559 425
rect -593 341 -559 357
rect -593 269 -559 289
rect -593 197 -559 221
rect -593 125 -559 153
rect -593 53 -559 85
rect -593 -17 -559 17
rect -593 -85 -559 -53
rect -593 -153 -559 -125
rect -593 -221 -559 -197
rect -593 -289 -559 -269
rect -593 -357 -559 -341
rect -593 -425 -559 -413
rect -593 -504 -559 -485
rect -497 485 -463 504
rect -497 413 -463 425
rect -497 341 -463 357
rect -497 269 -463 289
rect -497 197 -463 221
rect -497 125 -463 153
rect -497 53 -463 85
rect -497 -17 -463 17
rect -497 -85 -463 -53
rect -497 -153 -463 -125
rect -497 -221 -463 -197
rect -497 -289 -463 -269
rect -497 -357 -463 -341
rect -497 -425 -463 -413
rect -497 -504 -463 -485
rect -401 485 -367 504
rect -401 413 -367 425
rect -401 341 -367 357
rect -401 269 -367 289
rect -401 197 -367 221
rect -401 125 -367 153
rect -401 53 -367 85
rect -401 -17 -367 17
rect -401 -85 -367 -53
rect -401 -153 -367 -125
rect -401 -221 -367 -197
rect -401 -289 -367 -269
rect -401 -357 -367 -341
rect -401 -425 -367 -413
rect -401 -504 -367 -485
rect -305 485 -271 504
rect -305 413 -271 425
rect -305 341 -271 357
rect -305 269 -271 289
rect -305 197 -271 221
rect -305 125 -271 153
rect -305 53 -271 85
rect -305 -17 -271 17
rect -305 -85 -271 -53
rect -305 -153 -271 -125
rect -305 -221 -271 -197
rect -305 -289 -271 -269
rect -305 -357 -271 -341
rect -305 -425 -271 -413
rect -305 -504 -271 -485
rect -209 485 -175 504
rect -209 413 -175 425
rect -209 341 -175 357
rect -209 269 -175 289
rect -209 197 -175 221
rect -209 125 -175 153
rect -209 53 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -53
rect -209 -153 -175 -125
rect -209 -221 -175 -197
rect -209 -289 -175 -269
rect -209 -357 -175 -341
rect -209 -425 -175 -413
rect -209 -504 -175 -485
rect -113 485 -79 504
rect -113 413 -79 425
rect -113 341 -79 357
rect -113 269 -79 289
rect -113 197 -79 221
rect -113 125 -79 153
rect -113 53 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -53
rect -113 -153 -79 -125
rect -113 -221 -79 -197
rect -113 -289 -79 -269
rect -113 -357 -79 -341
rect -113 -425 -79 -413
rect -113 -504 -79 -485
rect -17 485 17 504
rect -17 413 17 425
rect -17 341 17 357
rect -17 269 17 289
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -289 17 -269
rect -17 -357 17 -341
rect -17 -425 17 -413
rect -17 -504 17 -485
rect 79 485 113 504
rect 79 413 113 425
rect 79 341 113 357
rect 79 269 113 289
rect 79 197 113 221
rect 79 125 113 153
rect 79 53 113 85
rect 79 -17 113 17
rect 79 -85 113 -53
rect 79 -153 113 -125
rect 79 -221 113 -197
rect 79 -289 113 -269
rect 79 -357 113 -341
rect 79 -425 113 -413
rect 79 -504 113 -485
rect 175 485 209 504
rect 175 413 209 425
rect 175 341 209 357
rect 175 269 209 289
rect 175 197 209 221
rect 175 125 209 153
rect 175 53 209 85
rect 175 -17 209 17
rect 175 -85 209 -53
rect 175 -153 209 -125
rect 175 -221 209 -197
rect 175 -289 209 -269
rect 175 -357 209 -341
rect 175 -425 209 -413
rect 175 -504 209 -485
rect 271 485 305 504
rect 271 413 305 425
rect 271 341 305 357
rect 271 269 305 289
rect 271 197 305 221
rect 271 125 305 153
rect 271 53 305 85
rect 271 -17 305 17
rect 271 -85 305 -53
rect 271 -153 305 -125
rect 271 -221 305 -197
rect 271 -289 305 -269
rect 271 -357 305 -341
rect 271 -425 305 -413
rect 271 -504 305 -485
rect 367 485 401 504
rect 367 413 401 425
rect 367 341 401 357
rect 367 269 401 289
rect 367 197 401 221
rect 367 125 401 153
rect 367 53 401 85
rect 367 -17 401 17
rect 367 -85 401 -53
rect 367 -153 401 -125
rect 367 -221 401 -197
rect 367 -289 401 -269
rect 367 -357 401 -341
rect 367 -425 401 -413
rect 367 -504 401 -485
rect 463 485 497 504
rect 463 413 497 425
rect 463 341 497 357
rect 463 269 497 289
rect 463 197 497 221
rect 463 125 497 153
rect 463 53 497 85
rect 463 -17 497 17
rect 463 -85 497 -53
rect 463 -153 497 -125
rect 463 -221 497 -197
rect 463 -289 497 -269
rect 463 -357 497 -341
rect 463 -425 497 -413
rect 463 -504 497 -485
rect 559 485 593 504
rect 559 413 593 425
rect 559 341 593 357
rect 559 269 593 289
rect 559 197 593 221
rect 559 125 593 153
rect 559 53 593 85
rect 559 -17 593 17
rect 559 -85 593 -53
rect 559 -153 593 -125
rect 559 -221 593 -197
rect 559 -289 593 -269
rect 559 -357 593 -341
rect 559 -425 593 -413
rect 559 -504 593 -485
rect 655 485 689 504
rect 655 413 689 425
rect 655 341 689 357
rect 655 269 689 289
rect 655 197 689 221
rect 655 125 689 153
rect 655 53 689 85
rect 655 -17 689 17
rect 655 -85 689 -53
rect 655 -153 689 -125
rect 655 -221 689 -197
rect 655 -289 689 -269
rect 655 -357 689 -341
rect 655 -425 689 -413
rect 655 -504 689 -485
rect 751 485 785 504
rect 751 413 785 425
rect 751 341 785 357
rect 751 269 785 289
rect 751 197 785 221
rect 751 125 785 153
rect 751 53 785 85
rect 751 -17 785 17
rect 751 -85 785 -53
rect 751 -153 785 -125
rect 751 -221 785 -197
rect 751 -289 785 -269
rect 751 -357 785 -341
rect 751 -425 785 -413
rect 751 -504 785 -485
rect 865 493 899 527
rect 865 425 899 459
rect 865 357 899 391
rect 865 289 899 323
rect 865 221 899 255
rect 865 153 899 187
rect 865 85 899 119
rect 865 17 899 51
rect 865 -51 899 -17
rect 865 -119 899 -85
rect 865 -187 899 -153
rect 865 -255 899 -221
rect 865 -323 899 -289
rect 865 -391 899 -357
rect 865 -459 899 -425
rect 865 -527 899 -493
rect -899 -649 -865 -561
rect -753 -581 -737 -547
rect -703 -581 -687 -547
rect -561 -581 -545 -547
rect -511 -581 -495 -547
rect -369 -581 -353 -547
rect -319 -581 -303 -547
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect 15 -581 31 -547
rect 65 -581 81 -547
rect 207 -581 223 -547
rect 257 -581 273 -547
rect 399 -581 415 -547
rect 449 -581 465 -547
rect 591 -581 607 -547
rect 641 -581 657 -547
rect 865 -649 899 -561
rect -899 -683 -799 -649
rect -765 -683 -731 -649
rect -697 -683 -663 -649
rect -629 -683 -595 -649
rect -561 -683 -527 -649
rect -493 -683 -459 -649
rect -425 -683 -391 -649
rect -357 -683 -323 -649
rect -289 -683 -255 -649
rect -221 -683 -187 -649
rect -153 -683 -119 -649
rect -85 -683 -51 -649
rect -17 -683 17 -649
rect 51 -683 85 -649
rect 119 -683 153 -649
rect 187 -683 221 -649
rect 255 -683 289 -649
rect 323 -683 357 -649
rect 391 -683 425 -649
rect 459 -683 493 -649
rect 527 -683 561 -649
rect 595 -683 629 -649
rect 663 -683 697 -649
rect 731 -683 765 -649
rect 799 -683 899 -649
<< viali >>
rect -641 547 -607 581
rect -449 547 -415 581
rect -257 547 -223 581
rect -65 547 -31 581
rect 127 547 161 581
rect 319 547 353 581
rect 511 547 545 581
rect 703 547 737 581
rect -785 459 -751 485
rect -785 451 -751 459
rect -785 391 -751 413
rect -785 379 -751 391
rect -785 323 -751 341
rect -785 307 -751 323
rect -785 255 -751 269
rect -785 235 -751 255
rect -785 187 -751 197
rect -785 163 -751 187
rect -785 119 -751 125
rect -785 91 -751 119
rect -785 51 -751 53
rect -785 19 -751 51
rect -785 -51 -751 -19
rect -785 -53 -751 -51
rect -785 -119 -751 -91
rect -785 -125 -751 -119
rect -785 -187 -751 -163
rect -785 -197 -751 -187
rect -785 -255 -751 -235
rect -785 -269 -751 -255
rect -785 -323 -751 -307
rect -785 -341 -751 -323
rect -785 -391 -751 -379
rect -785 -413 -751 -391
rect -785 -459 -751 -451
rect -785 -485 -751 -459
rect -689 459 -655 485
rect -689 451 -655 459
rect -689 391 -655 413
rect -689 379 -655 391
rect -689 323 -655 341
rect -689 307 -655 323
rect -689 255 -655 269
rect -689 235 -655 255
rect -689 187 -655 197
rect -689 163 -655 187
rect -689 119 -655 125
rect -689 91 -655 119
rect -689 51 -655 53
rect -689 19 -655 51
rect -689 -51 -655 -19
rect -689 -53 -655 -51
rect -689 -119 -655 -91
rect -689 -125 -655 -119
rect -689 -187 -655 -163
rect -689 -197 -655 -187
rect -689 -255 -655 -235
rect -689 -269 -655 -255
rect -689 -323 -655 -307
rect -689 -341 -655 -323
rect -689 -391 -655 -379
rect -689 -413 -655 -391
rect -689 -459 -655 -451
rect -689 -485 -655 -459
rect -593 459 -559 485
rect -593 451 -559 459
rect -593 391 -559 413
rect -593 379 -559 391
rect -593 323 -559 341
rect -593 307 -559 323
rect -593 255 -559 269
rect -593 235 -559 255
rect -593 187 -559 197
rect -593 163 -559 187
rect -593 119 -559 125
rect -593 91 -559 119
rect -593 51 -559 53
rect -593 19 -559 51
rect -593 -51 -559 -19
rect -593 -53 -559 -51
rect -593 -119 -559 -91
rect -593 -125 -559 -119
rect -593 -187 -559 -163
rect -593 -197 -559 -187
rect -593 -255 -559 -235
rect -593 -269 -559 -255
rect -593 -323 -559 -307
rect -593 -341 -559 -323
rect -593 -391 -559 -379
rect -593 -413 -559 -391
rect -593 -459 -559 -451
rect -593 -485 -559 -459
rect -497 459 -463 485
rect -497 451 -463 459
rect -497 391 -463 413
rect -497 379 -463 391
rect -497 323 -463 341
rect -497 307 -463 323
rect -497 255 -463 269
rect -497 235 -463 255
rect -497 187 -463 197
rect -497 163 -463 187
rect -497 119 -463 125
rect -497 91 -463 119
rect -497 51 -463 53
rect -497 19 -463 51
rect -497 -51 -463 -19
rect -497 -53 -463 -51
rect -497 -119 -463 -91
rect -497 -125 -463 -119
rect -497 -187 -463 -163
rect -497 -197 -463 -187
rect -497 -255 -463 -235
rect -497 -269 -463 -255
rect -497 -323 -463 -307
rect -497 -341 -463 -323
rect -497 -391 -463 -379
rect -497 -413 -463 -391
rect -497 -459 -463 -451
rect -497 -485 -463 -459
rect -401 459 -367 485
rect -401 451 -367 459
rect -401 391 -367 413
rect -401 379 -367 391
rect -401 323 -367 341
rect -401 307 -367 323
rect -401 255 -367 269
rect -401 235 -367 255
rect -401 187 -367 197
rect -401 163 -367 187
rect -401 119 -367 125
rect -401 91 -367 119
rect -401 51 -367 53
rect -401 19 -367 51
rect -401 -51 -367 -19
rect -401 -53 -367 -51
rect -401 -119 -367 -91
rect -401 -125 -367 -119
rect -401 -187 -367 -163
rect -401 -197 -367 -187
rect -401 -255 -367 -235
rect -401 -269 -367 -255
rect -401 -323 -367 -307
rect -401 -341 -367 -323
rect -401 -391 -367 -379
rect -401 -413 -367 -391
rect -401 -459 -367 -451
rect -401 -485 -367 -459
rect -305 459 -271 485
rect -305 451 -271 459
rect -305 391 -271 413
rect -305 379 -271 391
rect -305 323 -271 341
rect -305 307 -271 323
rect -305 255 -271 269
rect -305 235 -271 255
rect -305 187 -271 197
rect -305 163 -271 187
rect -305 119 -271 125
rect -305 91 -271 119
rect -305 51 -271 53
rect -305 19 -271 51
rect -305 -51 -271 -19
rect -305 -53 -271 -51
rect -305 -119 -271 -91
rect -305 -125 -271 -119
rect -305 -187 -271 -163
rect -305 -197 -271 -187
rect -305 -255 -271 -235
rect -305 -269 -271 -255
rect -305 -323 -271 -307
rect -305 -341 -271 -323
rect -305 -391 -271 -379
rect -305 -413 -271 -391
rect -305 -459 -271 -451
rect -305 -485 -271 -459
rect -209 459 -175 485
rect -209 451 -175 459
rect -209 391 -175 413
rect -209 379 -175 391
rect -209 323 -175 341
rect -209 307 -175 323
rect -209 255 -175 269
rect -209 235 -175 255
rect -209 187 -175 197
rect -209 163 -175 187
rect -209 119 -175 125
rect -209 91 -175 119
rect -209 51 -175 53
rect -209 19 -175 51
rect -209 -51 -175 -19
rect -209 -53 -175 -51
rect -209 -119 -175 -91
rect -209 -125 -175 -119
rect -209 -187 -175 -163
rect -209 -197 -175 -187
rect -209 -255 -175 -235
rect -209 -269 -175 -255
rect -209 -323 -175 -307
rect -209 -341 -175 -323
rect -209 -391 -175 -379
rect -209 -413 -175 -391
rect -209 -459 -175 -451
rect -209 -485 -175 -459
rect -113 459 -79 485
rect -113 451 -79 459
rect -113 391 -79 413
rect -113 379 -79 391
rect -113 323 -79 341
rect -113 307 -79 323
rect -113 255 -79 269
rect -113 235 -79 255
rect -113 187 -79 197
rect -113 163 -79 187
rect -113 119 -79 125
rect -113 91 -79 119
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -113 -119 -79 -91
rect -113 -125 -79 -119
rect -113 -187 -79 -163
rect -113 -197 -79 -187
rect -113 -255 -79 -235
rect -113 -269 -79 -255
rect -113 -323 -79 -307
rect -113 -341 -79 -323
rect -113 -391 -79 -379
rect -113 -413 -79 -391
rect -113 -459 -79 -451
rect -113 -485 -79 -459
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect 79 459 113 485
rect 79 451 113 459
rect 79 391 113 413
rect 79 379 113 391
rect 79 323 113 341
rect 79 307 113 323
rect 79 255 113 269
rect 79 235 113 255
rect 79 187 113 197
rect 79 163 113 187
rect 79 119 113 125
rect 79 91 113 119
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect 79 -119 113 -91
rect 79 -125 113 -119
rect 79 -187 113 -163
rect 79 -197 113 -187
rect 79 -255 113 -235
rect 79 -269 113 -255
rect 79 -323 113 -307
rect 79 -341 113 -323
rect 79 -391 113 -379
rect 79 -413 113 -391
rect 79 -459 113 -451
rect 79 -485 113 -459
rect 175 459 209 485
rect 175 451 209 459
rect 175 391 209 413
rect 175 379 209 391
rect 175 323 209 341
rect 175 307 209 323
rect 175 255 209 269
rect 175 235 209 255
rect 175 187 209 197
rect 175 163 209 187
rect 175 119 209 125
rect 175 91 209 119
rect 175 51 209 53
rect 175 19 209 51
rect 175 -51 209 -19
rect 175 -53 209 -51
rect 175 -119 209 -91
rect 175 -125 209 -119
rect 175 -187 209 -163
rect 175 -197 209 -187
rect 175 -255 209 -235
rect 175 -269 209 -255
rect 175 -323 209 -307
rect 175 -341 209 -323
rect 175 -391 209 -379
rect 175 -413 209 -391
rect 175 -459 209 -451
rect 175 -485 209 -459
rect 271 459 305 485
rect 271 451 305 459
rect 271 391 305 413
rect 271 379 305 391
rect 271 323 305 341
rect 271 307 305 323
rect 271 255 305 269
rect 271 235 305 255
rect 271 187 305 197
rect 271 163 305 187
rect 271 119 305 125
rect 271 91 305 119
rect 271 51 305 53
rect 271 19 305 51
rect 271 -51 305 -19
rect 271 -53 305 -51
rect 271 -119 305 -91
rect 271 -125 305 -119
rect 271 -187 305 -163
rect 271 -197 305 -187
rect 271 -255 305 -235
rect 271 -269 305 -255
rect 271 -323 305 -307
rect 271 -341 305 -323
rect 271 -391 305 -379
rect 271 -413 305 -391
rect 271 -459 305 -451
rect 271 -485 305 -459
rect 367 459 401 485
rect 367 451 401 459
rect 367 391 401 413
rect 367 379 401 391
rect 367 323 401 341
rect 367 307 401 323
rect 367 255 401 269
rect 367 235 401 255
rect 367 187 401 197
rect 367 163 401 187
rect 367 119 401 125
rect 367 91 401 119
rect 367 51 401 53
rect 367 19 401 51
rect 367 -51 401 -19
rect 367 -53 401 -51
rect 367 -119 401 -91
rect 367 -125 401 -119
rect 367 -187 401 -163
rect 367 -197 401 -187
rect 367 -255 401 -235
rect 367 -269 401 -255
rect 367 -323 401 -307
rect 367 -341 401 -323
rect 367 -391 401 -379
rect 367 -413 401 -391
rect 367 -459 401 -451
rect 367 -485 401 -459
rect 463 459 497 485
rect 463 451 497 459
rect 463 391 497 413
rect 463 379 497 391
rect 463 323 497 341
rect 463 307 497 323
rect 463 255 497 269
rect 463 235 497 255
rect 463 187 497 197
rect 463 163 497 187
rect 463 119 497 125
rect 463 91 497 119
rect 463 51 497 53
rect 463 19 497 51
rect 463 -51 497 -19
rect 463 -53 497 -51
rect 463 -119 497 -91
rect 463 -125 497 -119
rect 463 -187 497 -163
rect 463 -197 497 -187
rect 463 -255 497 -235
rect 463 -269 497 -255
rect 463 -323 497 -307
rect 463 -341 497 -323
rect 463 -391 497 -379
rect 463 -413 497 -391
rect 463 -459 497 -451
rect 463 -485 497 -459
rect 559 459 593 485
rect 559 451 593 459
rect 559 391 593 413
rect 559 379 593 391
rect 559 323 593 341
rect 559 307 593 323
rect 559 255 593 269
rect 559 235 593 255
rect 559 187 593 197
rect 559 163 593 187
rect 559 119 593 125
rect 559 91 593 119
rect 559 51 593 53
rect 559 19 593 51
rect 559 -51 593 -19
rect 559 -53 593 -51
rect 559 -119 593 -91
rect 559 -125 593 -119
rect 559 -187 593 -163
rect 559 -197 593 -187
rect 559 -255 593 -235
rect 559 -269 593 -255
rect 559 -323 593 -307
rect 559 -341 593 -323
rect 559 -391 593 -379
rect 559 -413 593 -391
rect 559 -459 593 -451
rect 559 -485 593 -459
rect 655 459 689 485
rect 655 451 689 459
rect 655 391 689 413
rect 655 379 689 391
rect 655 323 689 341
rect 655 307 689 323
rect 655 255 689 269
rect 655 235 689 255
rect 655 187 689 197
rect 655 163 689 187
rect 655 119 689 125
rect 655 91 689 119
rect 655 51 689 53
rect 655 19 689 51
rect 655 -51 689 -19
rect 655 -53 689 -51
rect 655 -119 689 -91
rect 655 -125 689 -119
rect 655 -187 689 -163
rect 655 -197 689 -187
rect 655 -255 689 -235
rect 655 -269 689 -255
rect 655 -323 689 -307
rect 655 -341 689 -323
rect 655 -391 689 -379
rect 655 -413 689 -391
rect 655 -459 689 -451
rect 655 -485 689 -459
rect 751 459 785 485
rect 751 451 785 459
rect 751 391 785 413
rect 751 379 785 391
rect 751 323 785 341
rect 751 307 785 323
rect 751 255 785 269
rect 751 235 785 255
rect 751 187 785 197
rect 751 163 785 187
rect 751 119 785 125
rect 751 91 785 119
rect 751 51 785 53
rect 751 19 785 51
rect 751 -51 785 -19
rect 751 -53 785 -51
rect 751 -119 785 -91
rect 751 -125 785 -119
rect 751 -187 785 -163
rect 751 -197 785 -187
rect 751 -255 785 -235
rect 751 -269 785 -255
rect 751 -323 785 -307
rect 751 -341 785 -323
rect 751 -391 785 -379
rect 751 -413 785 -391
rect 751 -459 785 -451
rect 751 -485 785 -459
rect -737 -581 -703 -547
rect -545 -581 -511 -547
rect -353 -581 -319 -547
rect -161 -581 -127 -547
rect 31 -581 65 -547
rect 223 -581 257 -547
rect 415 -581 449 -547
rect 607 -581 641 -547
<< metal1 >>
rect -653 581 -595 587
rect -653 547 -641 581
rect -607 547 -595 581
rect -653 541 -595 547
rect -461 581 -403 587
rect -461 547 -449 581
rect -415 547 -403 581
rect -461 541 -403 547
rect -269 581 -211 587
rect -269 547 -257 581
rect -223 547 -211 581
rect -269 541 -211 547
rect -77 581 -19 587
rect -77 547 -65 581
rect -31 547 -19 581
rect -77 541 -19 547
rect 115 581 173 587
rect 115 547 127 581
rect 161 547 173 581
rect 115 541 173 547
rect 307 581 365 587
rect 307 547 319 581
rect 353 547 365 581
rect 307 541 365 547
rect 499 581 557 587
rect 499 547 511 581
rect 545 547 557 581
rect 499 541 557 547
rect 691 581 749 587
rect 691 547 703 581
rect 737 547 749 581
rect 691 541 749 547
rect -791 485 -745 500
rect -791 451 -785 485
rect -751 451 -745 485
rect -791 413 -745 451
rect -791 379 -785 413
rect -751 379 -745 413
rect -791 341 -745 379
rect -791 307 -785 341
rect -751 307 -745 341
rect -791 269 -745 307
rect -791 235 -785 269
rect -751 235 -745 269
rect -791 197 -745 235
rect -791 163 -785 197
rect -751 163 -745 197
rect -791 125 -745 163
rect -791 91 -785 125
rect -751 91 -745 125
rect -791 53 -745 91
rect -791 19 -785 53
rect -751 19 -745 53
rect -791 -19 -745 19
rect -791 -53 -785 -19
rect -751 -53 -745 -19
rect -791 -91 -745 -53
rect -791 -125 -785 -91
rect -751 -125 -745 -91
rect -791 -163 -745 -125
rect -791 -197 -785 -163
rect -751 -197 -745 -163
rect -791 -235 -745 -197
rect -791 -269 -785 -235
rect -751 -269 -745 -235
rect -791 -307 -745 -269
rect -791 -341 -785 -307
rect -751 -341 -745 -307
rect -791 -379 -745 -341
rect -791 -413 -785 -379
rect -751 -413 -745 -379
rect -791 -451 -745 -413
rect -791 -485 -785 -451
rect -751 -485 -745 -451
rect -791 -500 -745 -485
rect -695 485 -649 500
rect -695 451 -689 485
rect -655 451 -649 485
rect -695 413 -649 451
rect -695 379 -689 413
rect -655 379 -649 413
rect -695 341 -649 379
rect -695 307 -689 341
rect -655 307 -649 341
rect -695 269 -649 307
rect -695 235 -689 269
rect -655 235 -649 269
rect -695 197 -649 235
rect -695 163 -689 197
rect -655 163 -649 197
rect -695 125 -649 163
rect -695 91 -689 125
rect -655 91 -649 125
rect -695 53 -649 91
rect -695 19 -689 53
rect -655 19 -649 53
rect -695 -19 -649 19
rect -695 -53 -689 -19
rect -655 -53 -649 -19
rect -695 -91 -649 -53
rect -695 -125 -689 -91
rect -655 -125 -649 -91
rect -695 -163 -649 -125
rect -695 -197 -689 -163
rect -655 -197 -649 -163
rect -695 -235 -649 -197
rect -695 -269 -689 -235
rect -655 -269 -649 -235
rect -695 -307 -649 -269
rect -695 -341 -689 -307
rect -655 -341 -649 -307
rect -695 -379 -649 -341
rect -695 -413 -689 -379
rect -655 -413 -649 -379
rect -695 -451 -649 -413
rect -695 -485 -689 -451
rect -655 -485 -649 -451
rect -695 -500 -649 -485
rect -599 485 -553 500
rect -599 451 -593 485
rect -559 451 -553 485
rect -599 413 -553 451
rect -599 379 -593 413
rect -559 379 -553 413
rect -599 341 -553 379
rect -599 307 -593 341
rect -559 307 -553 341
rect -599 269 -553 307
rect -599 235 -593 269
rect -559 235 -553 269
rect -599 197 -553 235
rect -599 163 -593 197
rect -559 163 -553 197
rect -599 125 -553 163
rect -599 91 -593 125
rect -559 91 -553 125
rect -599 53 -553 91
rect -599 19 -593 53
rect -559 19 -553 53
rect -599 -19 -553 19
rect -599 -53 -593 -19
rect -559 -53 -553 -19
rect -599 -91 -553 -53
rect -599 -125 -593 -91
rect -559 -125 -553 -91
rect -599 -163 -553 -125
rect -599 -197 -593 -163
rect -559 -197 -553 -163
rect -599 -235 -553 -197
rect -599 -269 -593 -235
rect -559 -269 -553 -235
rect -599 -307 -553 -269
rect -599 -341 -593 -307
rect -559 -341 -553 -307
rect -599 -379 -553 -341
rect -599 -413 -593 -379
rect -559 -413 -553 -379
rect -599 -451 -553 -413
rect -599 -485 -593 -451
rect -559 -485 -553 -451
rect -599 -500 -553 -485
rect -503 485 -457 500
rect -503 451 -497 485
rect -463 451 -457 485
rect -503 413 -457 451
rect -503 379 -497 413
rect -463 379 -457 413
rect -503 341 -457 379
rect -503 307 -497 341
rect -463 307 -457 341
rect -503 269 -457 307
rect -503 235 -497 269
rect -463 235 -457 269
rect -503 197 -457 235
rect -503 163 -497 197
rect -463 163 -457 197
rect -503 125 -457 163
rect -503 91 -497 125
rect -463 91 -457 125
rect -503 53 -457 91
rect -503 19 -497 53
rect -463 19 -457 53
rect -503 -19 -457 19
rect -503 -53 -497 -19
rect -463 -53 -457 -19
rect -503 -91 -457 -53
rect -503 -125 -497 -91
rect -463 -125 -457 -91
rect -503 -163 -457 -125
rect -503 -197 -497 -163
rect -463 -197 -457 -163
rect -503 -235 -457 -197
rect -503 -269 -497 -235
rect -463 -269 -457 -235
rect -503 -307 -457 -269
rect -503 -341 -497 -307
rect -463 -341 -457 -307
rect -503 -379 -457 -341
rect -503 -413 -497 -379
rect -463 -413 -457 -379
rect -503 -451 -457 -413
rect -503 -485 -497 -451
rect -463 -485 -457 -451
rect -503 -500 -457 -485
rect -407 485 -361 500
rect -407 451 -401 485
rect -367 451 -361 485
rect -407 413 -361 451
rect -407 379 -401 413
rect -367 379 -361 413
rect -407 341 -361 379
rect -407 307 -401 341
rect -367 307 -361 341
rect -407 269 -361 307
rect -407 235 -401 269
rect -367 235 -361 269
rect -407 197 -361 235
rect -407 163 -401 197
rect -367 163 -361 197
rect -407 125 -361 163
rect -407 91 -401 125
rect -367 91 -361 125
rect -407 53 -361 91
rect -407 19 -401 53
rect -367 19 -361 53
rect -407 -19 -361 19
rect -407 -53 -401 -19
rect -367 -53 -361 -19
rect -407 -91 -361 -53
rect -407 -125 -401 -91
rect -367 -125 -361 -91
rect -407 -163 -361 -125
rect -407 -197 -401 -163
rect -367 -197 -361 -163
rect -407 -235 -361 -197
rect -407 -269 -401 -235
rect -367 -269 -361 -235
rect -407 -307 -361 -269
rect -407 -341 -401 -307
rect -367 -341 -361 -307
rect -407 -379 -361 -341
rect -407 -413 -401 -379
rect -367 -413 -361 -379
rect -407 -451 -361 -413
rect -407 -485 -401 -451
rect -367 -485 -361 -451
rect -407 -500 -361 -485
rect -311 485 -265 500
rect -311 451 -305 485
rect -271 451 -265 485
rect -311 413 -265 451
rect -311 379 -305 413
rect -271 379 -265 413
rect -311 341 -265 379
rect -311 307 -305 341
rect -271 307 -265 341
rect -311 269 -265 307
rect -311 235 -305 269
rect -271 235 -265 269
rect -311 197 -265 235
rect -311 163 -305 197
rect -271 163 -265 197
rect -311 125 -265 163
rect -311 91 -305 125
rect -271 91 -265 125
rect -311 53 -265 91
rect -311 19 -305 53
rect -271 19 -265 53
rect -311 -19 -265 19
rect -311 -53 -305 -19
rect -271 -53 -265 -19
rect -311 -91 -265 -53
rect -311 -125 -305 -91
rect -271 -125 -265 -91
rect -311 -163 -265 -125
rect -311 -197 -305 -163
rect -271 -197 -265 -163
rect -311 -235 -265 -197
rect -311 -269 -305 -235
rect -271 -269 -265 -235
rect -311 -307 -265 -269
rect -311 -341 -305 -307
rect -271 -341 -265 -307
rect -311 -379 -265 -341
rect -311 -413 -305 -379
rect -271 -413 -265 -379
rect -311 -451 -265 -413
rect -311 -485 -305 -451
rect -271 -485 -265 -451
rect -311 -500 -265 -485
rect -215 485 -169 500
rect -215 451 -209 485
rect -175 451 -169 485
rect -215 413 -169 451
rect -215 379 -209 413
rect -175 379 -169 413
rect -215 341 -169 379
rect -215 307 -209 341
rect -175 307 -169 341
rect -215 269 -169 307
rect -215 235 -209 269
rect -175 235 -169 269
rect -215 197 -169 235
rect -215 163 -209 197
rect -175 163 -169 197
rect -215 125 -169 163
rect -215 91 -209 125
rect -175 91 -169 125
rect -215 53 -169 91
rect -215 19 -209 53
rect -175 19 -169 53
rect -215 -19 -169 19
rect -215 -53 -209 -19
rect -175 -53 -169 -19
rect -215 -91 -169 -53
rect -215 -125 -209 -91
rect -175 -125 -169 -91
rect -215 -163 -169 -125
rect -215 -197 -209 -163
rect -175 -197 -169 -163
rect -215 -235 -169 -197
rect -215 -269 -209 -235
rect -175 -269 -169 -235
rect -215 -307 -169 -269
rect -215 -341 -209 -307
rect -175 -341 -169 -307
rect -215 -379 -169 -341
rect -215 -413 -209 -379
rect -175 -413 -169 -379
rect -215 -451 -169 -413
rect -215 -485 -209 -451
rect -175 -485 -169 -451
rect -215 -500 -169 -485
rect -119 485 -73 500
rect -119 451 -113 485
rect -79 451 -73 485
rect -119 413 -73 451
rect -119 379 -113 413
rect -79 379 -73 413
rect -119 341 -73 379
rect -119 307 -113 341
rect -79 307 -73 341
rect -119 269 -73 307
rect -119 235 -113 269
rect -79 235 -73 269
rect -119 197 -73 235
rect -119 163 -113 197
rect -79 163 -73 197
rect -119 125 -73 163
rect -119 91 -113 125
rect -79 91 -73 125
rect -119 53 -73 91
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -91 -73 -53
rect -119 -125 -113 -91
rect -79 -125 -73 -91
rect -119 -163 -73 -125
rect -119 -197 -113 -163
rect -79 -197 -73 -163
rect -119 -235 -73 -197
rect -119 -269 -113 -235
rect -79 -269 -73 -235
rect -119 -307 -73 -269
rect -119 -341 -113 -307
rect -79 -341 -73 -307
rect -119 -379 -73 -341
rect -119 -413 -113 -379
rect -79 -413 -73 -379
rect -119 -451 -73 -413
rect -119 -485 -113 -451
rect -79 -485 -73 -451
rect -119 -500 -73 -485
rect -23 485 23 500
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -500 23 -485
rect 73 485 119 500
rect 73 451 79 485
rect 113 451 119 485
rect 73 413 119 451
rect 73 379 79 413
rect 113 379 119 413
rect 73 341 119 379
rect 73 307 79 341
rect 113 307 119 341
rect 73 269 119 307
rect 73 235 79 269
rect 113 235 119 269
rect 73 197 119 235
rect 73 163 79 197
rect 113 163 119 197
rect 73 125 119 163
rect 73 91 79 125
rect 113 91 119 125
rect 73 53 119 91
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -91 119 -53
rect 73 -125 79 -91
rect 113 -125 119 -91
rect 73 -163 119 -125
rect 73 -197 79 -163
rect 113 -197 119 -163
rect 73 -235 119 -197
rect 73 -269 79 -235
rect 113 -269 119 -235
rect 73 -307 119 -269
rect 73 -341 79 -307
rect 113 -341 119 -307
rect 73 -379 119 -341
rect 73 -413 79 -379
rect 113 -413 119 -379
rect 73 -451 119 -413
rect 73 -485 79 -451
rect 113 -485 119 -451
rect 73 -500 119 -485
rect 169 485 215 500
rect 169 451 175 485
rect 209 451 215 485
rect 169 413 215 451
rect 169 379 175 413
rect 209 379 215 413
rect 169 341 215 379
rect 169 307 175 341
rect 209 307 215 341
rect 169 269 215 307
rect 169 235 175 269
rect 209 235 215 269
rect 169 197 215 235
rect 169 163 175 197
rect 209 163 215 197
rect 169 125 215 163
rect 169 91 175 125
rect 209 91 215 125
rect 169 53 215 91
rect 169 19 175 53
rect 209 19 215 53
rect 169 -19 215 19
rect 169 -53 175 -19
rect 209 -53 215 -19
rect 169 -91 215 -53
rect 169 -125 175 -91
rect 209 -125 215 -91
rect 169 -163 215 -125
rect 169 -197 175 -163
rect 209 -197 215 -163
rect 169 -235 215 -197
rect 169 -269 175 -235
rect 209 -269 215 -235
rect 169 -307 215 -269
rect 169 -341 175 -307
rect 209 -341 215 -307
rect 169 -379 215 -341
rect 169 -413 175 -379
rect 209 -413 215 -379
rect 169 -451 215 -413
rect 169 -485 175 -451
rect 209 -485 215 -451
rect 169 -500 215 -485
rect 265 485 311 500
rect 265 451 271 485
rect 305 451 311 485
rect 265 413 311 451
rect 265 379 271 413
rect 305 379 311 413
rect 265 341 311 379
rect 265 307 271 341
rect 305 307 311 341
rect 265 269 311 307
rect 265 235 271 269
rect 305 235 311 269
rect 265 197 311 235
rect 265 163 271 197
rect 305 163 311 197
rect 265 125 311 163
rect 265 91 271 125
rect 305 91 311 125
rect 265 53 311 91
rect 265 19 271 53
rect 305 19 311 53
rect 265 -19 311 19
rect 265 -53 271 -19
rect 305 -53 311 -19
rect 265 -91 311 -53
rect 265 -125 271 -91
rect 305 -125 311 -91
rect 265 -163 311 -125
rect 265 -197 271 -163
rect 305 -197 311 -163
rect 265 -235 311 -197
rect 265 -269 271 -235
rect 305 -269 311 -235
rect 265 -307 311 -269
rect 265 -341 271 -307
rect 305 -341 311 -307
rect 265 -379 311 -341
rect 265 -413 271 -379
rect 305 -413 311 -379
rect 265 -451 311 -413
rect 265 -485 271 -451
rect 305 -485 311 -451
rect 265 -500 311 -485
rect 361 485 407 500
rect 361 451 367 485
rect 401 451 407 485
rect 361 413 407 451
rect 361 379 367 413
rect 401 379 407 413
rect 361 341 407 379
rect 361 307 367 341
rect 401 307 407 341
rect 361 269 407 307
rect 361 235 367 269
rect 401 235 407 269
rect 361 197 407 235
rect 361 163 367 197
rect 401 163 407 197
rect 361 125 407 163
rect 361 91 367 125
rect 401 91 407 125
rect 361 53 407 91
rect 361 19 367 53
rect 401 19 407 53
rect 361 -19 407 19
rect 361 -53 367 -19
rect 401 -53 407 -19
rect 361 -91 407 -53
rect 361 -125 367 -91
rect 401 -125 407 -91
rect 361 -163 407 -125
rect 361 -197 367 -163
rect 401 -197 407 -163
rect 361 -235 407 -197
rect 361 -269 367 -235
rect 401 -269 407 -235
rect 361 -307 407 -269
rect 361 -341 367 -307
rect 401 -341 407 -307
rect 361 -379 407 -341
rect 361 -413 367 -379
rect 401 -413 407 -379
rect 361 -451 407 -413
rect 361 -485 367 -451
rect 401 -485 407 -451
rect 361 -500 407 -485
rect 457 485 503 500
rect 457 451 463 485
rect 497 451 503 485
rect 457 413 503 451
rect 457 379 463 413
rect 497 379 503 413
rect 457 341 503 379
rect 457 307 463 341
rect 497 307 503 341
rect 457 269 503 307
rect 457 235 463 269
rect 497 235 503 269
rect 457 197 503 235
rect 457 163 463 197
rect 497 163 503 197
rect 457 125 503 163
rect 457 91 463 125
rect 497 91 503 125
rect 457 53 503 91
rect 457 19 463 53
rect 497 19 503 53
rect 457 -19 503 19
rect 457 -53 463 -19
rect 497 -53 503 -19
rect 457 -91 503 -53
rect 457 -125 463 -91
rect 497 -125 503 -91
rect 457 -163 503 -125
rect 457 -197 463 -163
rect 497 -197 503 -163
rect 457 -235 503 -197
rect 457 -269 463 -235
rect 497 -269 503 -235
rect 457 -307 503 -269
rect 457 -341 463 -307
rect 497 -341 503 -307
rect 457 -379 503 -341
rect 457 -413 463 -379
rect 497 -413 503 -379
rect 457 -451 503 -413
rect 457 -485 463 -451
rect 497 -485 503 -451
rect 457 -500 503 -485
rect 553 485 599 500
rect 553 451 559 485
rect 593 451 599 485
rect 553 413 599 451
rect 553 379 559 413
rect 593 379 599 413
rect 553 341 599 379
rect 553 307 559 341
rect 593 307 599 341
rect 553 269 599 307
rect 553 235 559 269
rect 593 235 599 269
rect 553 197 599 235
rect 553 163 559 197
rect 593 163 599 197
rect 553 125 599 163
rect 553 91 559 125
rect 593 91 599 125
rect 553 53 599 91
rect 553 19 559 53
rect 593 19 599 53
rect 553 -19 599 19
rect 553 -53 559 -19
rect 593 -53 599 -19
rect 553 -91 599 -53
rect 553 -125 559 -91
rect 593 -125 599 -91
rect 553 -163 599 -125
rect 553 -197 559 -163
rect 593 -197 599 -163
rect 553 -235 599 -197
rect 553 -269 559 -235
rect 593 -269 599 -235
rect 553 -307 599 -269
rect 553 -341 559 -307
rect 593 -341 599 -307
rect 553 -379 599 -341
rect 553 -413 559 -379
rect 593 -413 599 -379
rect 553 -451 599 -413
rect 553 -485 559 -451
rect 593 -485 599 -451
rect 553 -500 599 -485
rect 649 485 695 500
rect 649 451 655 485
rect 689 451 695 485
rect 649 413 695 451
rect 649 379 655 413
rect 689 379 695 413
rect 649 341 695 379
rect 649 307 655 341
rect 689 307 695 341
rect 649 269 695 307
rect 649 235 655 269
rect 689 235 695 269
rect 649 197 695 235
rect 649 163 655 197
rect 689 163 695 197
rect 649 125 695 163
rect 649 91 655 125
rect 689 91 695 125
rect 649 53 695 91
rect 649 19 655 53
rect 689 19 695 53
rect 649 -19 695 19
rect 649 -53 655 -19
rect 689 -53 695 -19
rect 649 -91 695 -53
rect 649 -125 655 -91
rect 689 -125 695 -91
rect 649 -163 695 -125
rect 649 -197 655 -163
rect 689 -197 695 -163
rect 649 -235 695 -197
rect 649 -269 655 -235
rect 689 -269 695 -235
rect 649 -307 695 -269
rect 649 -341 655 -307
rect 689 -341 695 -307
rect 649 -379 695 -341
rect 649 -413 655 -379
rect 689 -413 695 -379
rect 649 -451 695 -413
rect 649 -485 655 -451
rect 689 -485 695 -451
rect 649 -500 695 -485
rect 745 485 791 500
rect 745 451 751 485
rect 785 451 791 485
rect 745 413 791 451
rect 745 379 751 413
rect 785 379 791 413
rect 745 341 791 379
rect 745 307 751 341
rect 785 307 791 341
rect 745 269 791 307
rect 745 235 751 269
rect 785 235 791 269
rect 745 197 791 235
rect 745 163 751 197
rect 785 163 791 197
rect 745 125 791 163
rect 745 91 751 125
rect 785 91 791 125
rect 745 53 791 91
rect 745 19 751 53
rect 785 19 791 53
rect 745 -19 791 19
rect 745 -53 751 -19
rect 785 -53 791 -19
rect 745 -91 791 -53
rect 745 -125 751 -91
rect 785 -125 791 -91
rect 745 -163 791 -125
rect 745 -197 751 -163
rect 785 -197 791 -163
rect 745 -235 791 -197
rect 745 -269 751 -235
rect 785 -269 791 -235
rect 745 -307 791 -269
rect 745 -341 751 -307
rect 785 -341 791 -307
rect 745 -379 791 -341
rect 745 -413 751 -379
rect 785 -413 791 -379
rect 745 -451 791 -413
rect 745 -485 751 -451
rect 785 -485 791 -451
rect 745 -500 791 -485
rect -749 -547 -691 -541
rect -749 -581 -737 -547
rect -703 -581 -691 -547
rect -749 -587 -691 -581
rect -557 -547 -499 -541
rect -557 -581 -545 -547
rect -511 -581 -499 -547
rect -557 -587 -499 -581
rect -365 -547 -307 -541
rect -365 -581 -353 -547
rect -319 -581 -307 -547
rect -365 -587 -307 -581
rect -173 -547 -115 -541
rect -173 -581 -161 -547
rect -127 -581 -115 -547
rect -173 -587 -115 -581
rect 19 -547 77 -541
rect 19 -581 31 -547
rect 65 -581 77 -547
rect 19 -587 77 -581
rect 211 -547 269 -541
rect 211 -581 223 -547
rect 257 -581 269 -547
rect 211 -587 269 -581
rect 403 -547 461 -541
rect 403 -581 415 -547
rect 449 -581 461 -547
rect 403 -587 461 -581
rect 595 -547 653 -541
rect 595 -581 607 -547
rect 641 -581 653 -547
rect 595 -587 653 -581
<< properties >>
string FIXED_BBOX -882 -666 882 666
<< end >>
