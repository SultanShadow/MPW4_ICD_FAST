magic
tech sky130A
magscale 1 2
timestamp 1640969486
<< poly >>
rect 56 539 5287 578
rect 56 505 86 539
rect 120 505 154 539
rect 188 505 222 539
rect 256 505 290 539
rect 324 505 358 539
rect 392 505 426 539
rect 460 505 494 539
rect 528 505 562 539
rect 596 505 630 539
rect 664 505 698 539
rect 732 505 766 539
rect 800 505 834 539
rect 868 505 902 539
rect 936 505 970 539
rect 1004 505 1038 539
rect 1072 505 1106 539
rect 1140 505 1174 539
rect 1208 505 1242 539
rect 1276 505 1310 539
rect 1344 505 1378 539
rect 1412 505 1446 539
rect 1480 505 1514 539
rect 1548 505 1582 539
rect 1616 505 1650 539
rect 1684 505 1718 539
rect 1752 505 1786 539
rect 1820 505 1854 539
rect 1888 505 1922 539
rect 1956 505 1990 539
rect 2024 505 2058 539
rect 2092 505 2126 539
rect 2160 505 2194 539
rect 2228 505 2262 539
rect 2296 505 2330 539
rect 2364 505 2398 539
rect 2432 505 2466 539
rect 2500 505 2534 539
rect 2568 505 2602 539
rect 2636 505 2670 539
rect 2704 505 2738 539
rect 2772 505 2806 539
rect 2840 505 2874 539
rect 2908 505 2942 539
rect 2976 505 3010 539
rect 3044 505 3078 539
rect 3112 505 3146 539
rect 3180 505 3214 539
rect 3248 505 3282 539
rect 3316 505 3350 539
rect 3384 505 3418 539
rect 3452 505 3486 539
rect 3520 505 3554 539
rect 3588 505 3622 539
rect 3656 505 3690 539
rect 3724 505 3758 539
rect 3792 505 3826 539
rect 3860 505 3894 539
rect 3928 505 3962 539
rect 3996 505 4030 539
rect 4064 505 4098 539
rect 4132 505 4166 539
rect 4200 505 4234 539
rect 4268 505 4302 539
rect 4336 505 4370 539
rect 4404 505 4438 539
rect 4472 505 4506 539
rect 4540 505 4574 539
rect 4608 505 4642 539
rect 4676 505 4710 539
rect 4744 505 4778 539
rect 4812 505 4846 539
rect 4880 505 4914 539
rect 4948 505 4982 539
rect 5016 505 5050 539
rect 5084 505 5118 539
rect 5152 505 5186 539
rect 5220 505 5287 539
rect 56 488 5287 505
rect 56 483 5288 488
rect 56 452 1056 483
rect 1114 452 2114 483
rect 2172 452 3172 483
rect 3230 452 4230 483
rect 4288 452 5288 483
<< polycont >>
rect 86 505 120 539
rect 154 505 188 539
rect 222 505 256 539
rect 290 505 324 539
rect 358 505 392 539
rect 426 505 460 539
rect 494 505 528 539
rect 562 505 596 539
rect 630 505 664 539
rect 698 505 732 539
rect 766 505 800 539
rect 834 505 868 539
rect 902 505 936 539
rect 970 505 1004 539
rect 1038 505 1072 539
rect 1106 505 1140 539
rect 1174 505 1208 539
rect 1242 505 1276 539
rect 1310 505 1344 539
rect 1378 505 1412 539
rect 1446 505 1480 539
rect 1514 505 1548 539
rect 1582 505 1616 539
rect 1650 505 1684 539
rect 1718 505 1752 539
rect 1786 505 1820 539
rect 1854 505 1888 539
rect 1922 505 1956 539
rect 1990 505 2024 539
rect 2058 505 2092 539
rect 2126 505 2160 539
rect 2194 505 2228 539
rect 2262 505 2296 539
rect 2330 505 2364 539
rect 2398 505 2432 539
rect 2466 505 2500 539
rect 2534 505 2568 539
rect 2602 505 2636 539
rect 2670 505 2704 539
rect 2738 505 2772 539
rect 2806 505 2840 539
rect 2874 505 2908 539
rect 2942 505 2976 539
rect 3010 505 3044 539
rect 3078 505 3112 539
rect 3146 505 3180 539
rect 3214 505 3248 539
rect 3282 505 3316 539
rect 3350 505 3384 539
rect 3418 505 3452 539
rect 3486 505 3520 539
rect 3554 505 3588 539
rect 3622 505 3656 539
rect 3690 505 3724 539
rect 3758 505 3792 539
rect 3826 505 3860 539
rect 3894 505 3928 539
rect 3962 505 3996 539
rect 4030 505 4064 539
rect 4098 505 4132 539
rect 4166 505 4200 539
rect 4234 505 4268 539
rect 4302 505 4336 539
rect 4370 505 4404 539
rect 4438 505 4472 539
rect 4506 505 4540 539
rect 4574 505 4608 539
rect 4642 505 4676 539
rect 4710 505 4744 539
rect 4778 505 4812 539
rect 4846 505 4880 539
rect 4914 505 4948 539
rect 4982 505 5016 539
rect 5050 505 5084 539
rect 5118 505 5152 539
rect 5186 505 5220 539
<< locali >>
rect 56 542 5287 578
rect 56 508 80 542
rect 114 539 152 542
rect 186 539 224 542
rect 258 539 296 542
rect 330 539 368 542
rect 402 539 440 542
rect 474 539 512 542
rect 546 539 584 542
rect 618 539 656 542
rect 690 539 728 542
rect 762 539 800 542
rect 120 508 152 539
rect 56 505 86 508
rect 120 505 154 508
rect 188 505 222 539
rect 258 508 290 539
rect 330 508 358 539
rect 402 508 426 539
rect 474 508 494 539
rect 546 508 562 539
rect 618 508 630 539
rect 690 508 698 539
rect 762 508 766 539
rect 256 505 290 508
rect 324 505 358 508
rect 392 505 426 508
rect 460 505 494 508
rect 528 505 562 508
rect 596 505 630 508
rect 664 505 698 508
rect 732 505 766 508
rect 834 539 872 542
rect 906 539 944 542
rect 978 539 1016 542
rect 1050 539 1088 542
rect 1122 539 1160 542
rect 1194 539 1232 542
rect 1266 539 1304 542
rect 1338 539 1376 542
rect 1410 539 1448 542
rect 1482 539 1520 542
rect 1554 539 1592 542
rect 1626 539 1664 542
rect 1698 539 1736 542
rect 1770 539 1808 542
rect 1842 539 1880 542
rect 1914 539 1952 542
rect 1986 539 2024 542
rect 800 505 834 508
rect 868 508 872 539
rect 936 508 944 539
rect 1004 508 1016 539
rect 1072 508 1088 539
rect 1140 508 1160 539
rect 1208 508 1232 539
rect 1276 508 1304 539
rect 1344 508 1376 539
rect 868 505 902 508
rect 936 505 970 508
rect 1004 505 1038 508
rect 1072 505 1106 508
rect 1140 505 1174 508
rect 1208 505 1242 508
rect 1276 505 1310 508
rect 1344 505 1378 508
rect 1412 505 1446 539
rect 1482 508 1514 539
rect 1554 508 1582 539
rect 1626 508 1650 539
rect 1698 508 1718 539
rect 1770 508 1786 539
rect 1842 508 1854 539
rect 1914 508 1922 539
rect 1986 508 1990 539
rect 1480 505 1514 508
rect 1548 505 1582 508
rect 1616 505 1650 508
rect 1684 505 1718 508
rect 1752 505 1786 508
rect 1820 505 1854 508
rect 1888 505 1922 508
rect 1956 505 1990 508
rect 2058 539 2096 542
rect 2130 539 2168 542
rect 2202 539 2240 542
rect 2274 539 2312 542
rect 2346 539 2384 542
rect 2418 539 2456 542
rect 2490 539 2528 542
rect 2562 539 2600 542
rect 2634 539 2672 542
rect 2706 539 2744 542
rect 2778 539 2816 542
rect 2850 539 2888 542
rect 2922 539 2960 542
rect 2994 539 3032 542
rect 3066 539 3104 542
rect 3138 539 3176 542
rect 3210 539 3248 542
rect 2024 505 2058 508
rect 2092 508 2096 539
rect 2160 508 2168 539
rect 2228 508 2240 539
rect 2296 508 2312 539
rect 2364 508 2384 539
rect 2432 508 2456 539
rect 2500 508 2528 539
rect 2568 508 2600 539
rect 2092 505 2126 508
rect 2160 505 2194 508
rect 2228 505 2262 508
rect 2296 505 2330 508
rect 2364 505 2398 508
rect 2432 505 2466 508
rect 2500 505 2534 508
rect 2568 505 2602 508
rect 2636 505 2670 539
rect 2706 508 2738 539
rect 2778 508 2806 539
rect 2850 508 2874 539
rect 2922 508 2942 539
rect 2994 508 3010 539
rect 3066 508 3078 539
rect 3138 508 3146 539
rect 3210 508 3214 539
rect 2704 505 2738 508
rect 2772 505 2806 508
rect 2840 505 2874 508
rect 2908 505 2942 508
rect 2976 505 3010 508
rect 3044 505 3078 508
rect 3112 505 3146 508
rect 3180 505 3214 508
rect 3282 539 3320 542
rect 3354 539 3392 542
rect 3426 539 3464 542
rect 3498 539 3536 542
rect 3570 539 3608 542
rect 3642 539 3680 542
rect 3714 539 3752 542
rect 3786 539 3824 542
rect 3858 539 3896 542
rect 3930 539 3968 542
rect 4002 539 4040 542
rect 4074 539 4112 542
rect 4146 539 4184 542
rect 4218 539 4256 542
rect 4290 539 4328 542
rect 4362 539 4400 542
rect 4434 539 4472 542
rect 3248 505 3282 508
rect 3316 508 3320 539
rect 3384 508 3392 539
rect 3452 508 3464 539
rect 3520 508 3536 539
rect 3588 508 3608 539
rect 3656 508 3680 539
rect 3724 508 3752 539
rect 3792 508 3824 539
rect 3316 505 3350 508
rect 3384 505 3418 508
rect 3452 505 3486 508
rect 3520 505 3554 508
rect 3588 505 3622 508
rect 3656 505 3690 508
rect 3724 505 3758 508
rect 3792 505 3826 508
rect 3860 505 3894 539
rect 3930 508 3962 539
rect 4002 508 4030 539
rect 4074 508 4098 539
rect 4146 508 4166 539
rect 4218 508 4234 539
rect 4290 508 4302 539
rect 4362 508 4370 539
rect 4434 508 4438 539
rect 3928 505 3962 508
rect 3996 505 4030 508
rect 4064 505 4098 508
rect 4132 505 4166 508
rect 4200 505 4234 508
rect 4268 505 4302 508
rect 4336 505 4370 508
rect 4404 505 4438 508
rect 4506 539 4544 542
rect 4578 539 4616 542
rect 4650 539 4688 542
rect 4722 539 4760 542
rect 4794 539 4832 542
rect 4866 539 4904 542
rect 4938 539 4976 542
rect 5010 539 5048 542
rect 5082 539 5120 542
rect 5154 539 5192 542
rect 4472 505 4506 508
rect 4540 508 4544 539
rect 4608 508 4616 539
rect 4676 508 4688 539
rect 4744 508 4760 539
rect 4812 508 4832 539
rect 4880 508 4904 539
rect 4948 508 4976 539
rect 5016 508 5048 539
rect 4540 505 4574 508
rect 4608 505 4642 508
rect 4676 505 4710 508
rect 4744 505 4778 508
rect 4812 505 4846 508
rect 4880 505 4914 508
rect 4948 505 4982 508
rect 5016 505 5050 508
rect 5084 505 5118 539
rect 5154 508 5186 539
rect 5226 508 5287 542
rect 5152 505 5186 508
rect 5220 505 5287 508
rect 56 483 5287 505
rect 1068 -20 1102 26
rect 3184 -20 3218 26
rect 5300 -20 5334 26
rect 1068 -102 5336 -20
<< viali >>
rect 80 539 114 542
rect 152 539 186 542
rect 224 539 258 542
rect 296 539 330 542
rect 368 539 402 542
rect 440 539 474 542
rect 512 539 546 542
rect 584 539 618 542
rect 656 539 690 542
rect 728 539 762 542
rect 80 508 86 539
rect 86 508 114 539
rect 152 508 154 539
rect 154 508 186 539
rect 224 508 256 539
rect 256 508 258 539
rect 296 508 324 539
rect 324 508 330 539
rect 368 508 392 539
rect 392 508 402 539
rect 440 508 460 539
rect 460 508 474 539
rect 512 508 528 539
rect 528 508 546 539
rect 584 508 596 539
rect 596 508 618 539
rect 656 508 664 539
rect 664 508 690 539
rect 728 508 732 539
rect 732 508 762 539
rect 800 508 834 542
rect 872 539 906 542
rect 944 539 978 542
rect 1016 539 1050 542
rect 1088 539 1122 542
rect 1160 539 1194 542
rect 1232 539 1266 542
rect 1304 539 1338 542
rect 1376 539 1410 542
rect 1448 539 1482 542
rect 1520 539 1554 542
rect 1592 539 1626 542
rect 1664 539 1698 542
rect 1736 539 1770 542
rect 1808 539 1842 542
rect 1880 539 1914 542
rect 1952 539 1986 542
rect 872 508 902 539
rect 902 508 906 539
rect 944 508 970 539
rect 970 508 978 539
rect 1016 508 1038 539
rect 1038 508 1050 539
rect 1088 508 1106 539
rect 1106 508 1122 539
rect 1160 508 1174 539
rect 1174 508 1194 539
rect 1232 508 1242 539
rect 1242 508 1266 539
rect 1304 508 1310 539
rect 1310 508 1338 539
rect 1376 508 1378 539
rect 1378 508 1410 539
rect 1448 508 1480 539
rect 1480 508 1482 539
rect 1520 508 1548 539
rect 1548 508 1554 539
rect 1592 508 1616 539
rect 1616 508 1626 539
rect 1664 508 1684 539
rect 1684 508 1698 539
rect 1736 508 1752 539
rect 1752 508 1770 539
rect 1808 508 1820 539
rect 1820 508 1842 539
rect 1880 508 1888 539
rect 1888 508 1914 539
rect 1952 508 1956 539
rect 1956 508 1986 539
rect 2024 508 2058 542
rect 2096 539 2130 542
rect 2168 539 2202 542
rect 2240 539 2274 542
rect 2312 539 2346 542
rect 2384 539 2418 542
rect 2456 539 2490 542
rect 2528 539 2562 542
rect 2600 539 2634 542
rect 2672 539 2706 542
rect 2744 539 2778 542
rect 2816 539 2850 542
rect 2888 539 2922 542
rect 2960 539 2994 542
rect 3032 539 3066 542
rect 3104 539 3138 542
rect 3176 539 3210 542
rect 2096 508 2126 539
rect 2126 508 2130 539
rect 2168 508 2194 539
rect 2194 508 2202 539
rect 2240 508 2262 539
rect 2262 508 2274 539
rect 2312 508 2330 539
rect 2330 508 2346 539
rect 2384 508 2398 539
rect 2398 508 2418 539
rect 2456 508 2466 539
rect 2466 508 2490 539
rect 2528 508 2534 539
rect 2534 508 2562 539
rect 2600 508 2602 539
rect 2602 508 2634 539
rect 2672 508 2704 539
rect 2704 508 2706 539
rect 2744 508 2772 539
rect 2772 508 2778 539
rect 2816 508 2840 539
rect 2840 508 2850 539
rect 2888 508 2908 539
rect 2908 508 2922 539
rect 2960 508 2976 539
rect 2976 508 2994 539
rect 3032 508 3044 539
rect 3044 508 3066 539
rect 3104 508 3112 539
rect 3112 508 3138 539
rect 3176 508 3180 539
rect 3180 508 3210 539
rect 3248 508 3282 542
rect 3320 539 3354 542
rect 3392 539 3426 542
rect 3464 539 3498 542
rect 3536 539 3570 542
rect 3608 539 3642 542
rect 3680 539 3714 542
rect 3752 539 3786 542
rect 3824 539 3858 542
rect 3896 539 3930 542
rect 3968 539 4002 542
rect 4040 539 4074 542
rect 4112 539 4146 542
rect 4184 539 4218 542
rect 4256 539 4290 542
rect 4328 539 4362 542
rect 4400 539 4434 542
rect 3320 508 3350 539
rect 3350 508 3354 539
rect 3392 508 3418 539
rect 3418 508 3426 539
rect 3464 508 3486 539
rect 3486 508 3498 539
rect 3536 508 3554 539
rect 3554 508 3570 539
rect 3608 508 3622 539
rect 3622 508 3642 539
rect 3680 508 3690 539
rect 3690 508 3714 539
rect 3752 508 3758 539
rect 3758 508 3786 539
rect 3824 508 3826 539
rect 3826 508 3858 539
rect 3896 508 3928 539
rect 3928 508 3930 539
rect 3968 508 3996 539
rect 3996 508 4002 539
rect 4040 508 4064 539
rect 4064 508 4074 539
rect 4112 508 4132 539
rect 4132 508 4146 539
rect 4184 508 4200 539
rect 4200 508 4218 539
rect 4256 508 4268 539
rect 4268 508 4290 539
rect 4328 508 4336 539
rect 4336 508 4362 539
rect 4400 508 4404 539
rect 4404 508 4434 539
rect 4472 508 4506 542
rect 4544 539 4578 542
rect 4616 539 4650 542
rect 4688 539 4722 542
rect 4760 539 4794 542
rect 4832 539 4866 542
rect 4904 539 4938 542
rect 4976 539 5010 542
rect 5048 539 5082 542
rect 5120 539 5154 542
rect 5192 539 5226 542
rect 4544 508 4574 539
rect 4574 508 4578 539
rect 4616 508 4642 539
rect 4642 508 4650 539
rect 4688 508 4710 539
rect 4710 508 4722 539
rect 4760 508 4778 539
rect 4778 508 4794 539
rect 4832 508 4846 539
rect 4846 508 4866 539
rect 4904 508 4914 539
rect 4914 508 4938 539
rect 4976 508 4982 539
rect 4982 508 5010 539
rect 5048 508 5050 539
rect 5050 508 5082 539
rect 5120 508 5152 539
rect 5152 508 5154 539
rect 5192 508 5220 539
rect 5220 508 5226 539
<< metal1 >>
rect 56 542 5288 578
rect 56 508 80 542
rect 114 508 152 542
rect 186 508 224 542
rect 258 508 296 542
rect 330 508 368 542
rect 402 508 440 542
rect 474 508 512 542
rect 546 508 584 542
rect 618 508 656 542
rect 690 508 728 542
rect 762 508 800 542
rect 834 508 872 542
rect 906 508 944 542
rect 978 508 1016 542
rect 1050 508 1088 542
rect 1122 508 1160 542
rect 1194 508 1232 542
rect 1266 508 1304 542
rect 1338 508 1376 542
rect 1410 508 1448 542
rect 1482 508 1520 542
rect 1554 508 1592 542
rect 1626 508 1664 542
rect 1698 508 1736 542
rect 1770 508 1808 542
rect 1842 508 1880 542
rect 1914 508 1952 542
rect 1986 508 2024 542
rect 2058 508 2096 542
rect 2130 508 2168 542
rect 2202 508 2240 542
rect 2274 508 2312 542
rect 2346 508 2384 542
rect 2418 508 2456 542
rect 2490 508 2528 542
rect 2562 508 2600 542
rect 2634 508 2672 542
rect 2706 508 2744 542
rect 2778 508 2816 542
rect 2850 508 2888 542
rect 2922 508 2960 542
rect 2994 508 3032 542
rect 3066 508 3104 542
rect 3138 508 3176 542
rect 3210 508 3248 542
rect 3282 508 3320 542
rect 3354 508 3392 542
rect 3426 508 3464 542
rect 3498 508 3536 542
rect 3570 508 3608 542
rect 3642 508 3680 542
rect 3714 508 3752 542
rect 3786 508 3824 542
rect 3858 508 3896 542
rect 3930 508 3968 542
rect 4002 508 4040 542
rect 4074 508 4112 542
rect 4146 508 4184 542
rect 4218 508 4256 542
rect 4290 508 4328 542
rect 4362 508 4400 542
rect 4434 508 4472 542
rect 4506 508 4544 542
rect 4578 508 4616 542
rect 4650 508 4688 542
rect 4722 508 4760 542
rect 4794 508 4832 542
rect 4866 508 4904 542
rect 4938 508 4976 542
rect 5010 508 5048 542
rect 5082 508 5120 542
rect 5154 508 5192 542
rect 5226 508 5288 542
rect 56 483 5288 508
rect 4 -21 50 28
rect 2120 -21 2166 28
rect 4236 -21 4282 28
rect 3 -123 4282 -21
use sky130_fd_pr__nfet_g5v0d10v5_CPNAJY  sky130_fd_pr__nfet_g5v0d10v5_CPNAJY_0
timestamp 1640969486
transform 1 0 556 0 1 226
box -584 -226 584 226
use sky130_fd_pr__nfet_g5v0d10v5_CPNAJY  sky130_fd_pr__nfet_g5v0d10v5_CPNAJY_1
timestamp 1640969486
transform 1 0 1614 0 1 226
box -584 -226 584 226
use sky130_fd_pr__nfet_g5v0d10v5_CPNAJY  sky130_fd_pr__nfet_g5v0d10v5_CPNAJY_2
timestamp 1640969486
transform 1 0 2672 0 1 226
box -584 -226 584 226
use sky130_fd_pr__nfet_g5v0d10v5_CPNAJY  sky130_fd_pr__nfet_g5v0d10v5_CPNAJY_3
timestamp 1640969486
transform 1 0 3730 0 1 226
box -584 -226 584 226
use sky130_fd_pr__nfet_g5v0d10v5_CPNAJY  sky130_fd_pr__nfet_g5v0d10v5_CPNAJY_4
timestamp 1640969486
transform 1 0 4788 0 1 226
box -584 -226 584 226
<< labels >>
flabel metal1 s 2426 558 2426 558 0 FreeSans 250 0 0 0 G
port 1 nsew
flabel metal1 s 300 -75 300 -75 0 FreeSans 250 0 0 0 D
port 2 nsew
flabel locali s 4646 -77 4646 -77 0 FreeSans 250 0 0 0 S
port 3 nsew
<< end >>
