magic
tech sky130A
magscale 1 2
timestamp 1640969486
<< error_p >>
rect -624 262 624 266
rect -624 -262 -594 262
rect -558 196 558 200
rect -558 -196 -528 196
rect 528 -196 558 196
rect -558 -200 558 -196
rect 594 -262 624 262
rect -624 -266 624 -262
<< nwell >>
rect -594 -262 594 262
<< mvpmos >>
rect -500 -200 500 200
<< mvpdiff >>
rect -558 187 -500 200
rect -558 153 -546 187
rect -512 153 -500 187
rect -558 119 -500 153
rect -558 85 -546 119
rect -512 85 -500 119
rect -558 51 -500 85
rect -558 17 -546 51
rect -512 17 -500 51
rect -558 -17 -500 17
rect -558 -51 -546 -17
rect -512 -51 -500 -17
rect -558 -85 -500 -51
rect -558 -119 -546 -85
rect -512 -119 -500 -85
rect -558 -153 -500 -119
rect -558 -187 -546 -153
rect -512 -187 -500 -153
rect -558 -200 -500 -187
rect 500 187 558 200
rect 500 153 512 187
rect 546 153 558 187
rect 500 119 558 153
rect 500 85 512 119
rect 546 85 558 119
rect 500 51 558 85
rect 500 17 512 51
rect 546 17 558 51
rect 500 -17 558 17
rect 500 -51 512 -17
rect 546 -51 558 -17
rect 500 -85 558 -51
rect 500 -119 512 -85
rect 546 -119 558 -85
rect 500 -153 558 -119
rect 500 -187 512 -153
rect 546 -187 558 -153
rect 500 -200 558 -187
<< mvpdiffc >>
rect -546 153 -512 187
rect -546 85 -512 119
rect -546 17 -512 51
rect -546 -51 -512 -17
rect -546 -119 -512 -85
rect -546 -187 -512 -153
rect 512 153 546 187
rect 512 85 546 119
rect 512 17 546 51
rect 512 -51 546 -17
rect 512 -119 546 -85
rect 512 -187 546 -153
<< poly >>
rect -500 200 500 226
rect -500 -226 500 -200
<< locali >>
rect -546 187 -512 204
rect -546 119 -512 127
rect -546 51 -512 55
rect -546 -55 -512 -51
rect -546 -127 -512 -119
rect -546 -204 -512 -187
rect 512 187 546 204
rect 512 119 546 127
rect 512 51 546 55
rect 512 -55 546 -51
rect 512 -127 546 -119
rect 512 -204 546 -187
<< viali >>
rect -546 153 -512 161
rect -546 127 -512 153
rect -546 85 -512 89
rect -546 55 -512 85
rect -546 -17 -512 17
rect -546 -85 -512 -55
rect -546 -89 -512 -85
rect -546 -153 -512 -127
rect -546 -161 -512 -153
rect 512 153 546 161
rect 512 127 546 153
rect 512 85 546 89
rect 512 55 546 85
rect 512 -17 546 17
rect 512 -85 546 -55
rect 512 -89 546 -85
rect 512 -153 546 -127
rect 512 -161 546 -153
<< metal1 >>
rect -552 161 -506 200
rect -552 127 -546 161
rect -512 127 -506 161
rect -552 89 -506 127
rect -552 55 -546 89
rect -512 55 -506 89
rect -552 17 -506 55
rect -552 -17 -546 17
rect -512 -17 -506 17
rect -552 -55 -506 -17
rect -552 -89 -546 -55
rect -512 -89 -506 -55
rect -552 -127 -506 -89
rect -552 -161 -546 -127
rect -512 -161 -506 -127
rect -552 -200 -506 -161
rect 506 161 552 200
rect 506 127 512 161
rect 546 127 552 161
rect 506 89 552 127
rect 506 55 512 89
rect 546 55 552 89
rect 506 17 552 55
rect 506 -17 512 17
rect 546 -17 552 17
rect 506 -55 552 -17
rect 506 -89 512 -55
rect 546 -89 552 -55
rect 506 -127 552 -89
rect 506 -161 512 -127
rect 546 -161 552 -127
rect 506 -200 552 -161
<< end >>
