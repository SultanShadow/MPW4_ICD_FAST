magic
tech sky130A
timestamp 1640969486
use FINAL_without_ind  FINAL_without_ind_0
timestamp 1640969486
transform 1 0 3570 0 1 0
box -3578 0 68406 49393
<< end >>
