magic
tech sky130A
magscale 1 2
timestamp 1640969486
<< nwell >>
rect -508 -541 3769 1749
<< nsubdiff >>
rect -347 1672 3631 1678
rect -347 1502 152 1672
rect 3178 1502 3631 1672
rect -347 1497 3631 1502
rect -347 1260 -129 1497
rect 3413 1312 3631 1497
rect -347 2 -323 1260
rect -153 2 -129 1260
rect 3413 54 3437 1312
rect 3607 54 3631 1312
rect -347 -184 -129 2
rect 3413 -184 3631 54
rect -347 -190 3631 -184
rect -347 -360 248 -190
rect 3274 -360 3631 -190
rect -347 -365 3631 -360
<< nsubdiffcont >>
rect 152 1502 3178 1672
rect -323 2 -153 1260
rect 3437 54 3607 1312
rect 248 -360 3274 -190
<< poly >>
rect 94 1380 3196 1394
rect 94 1346 123 1380
rect 157 1346 191 1380
rect 225 1346 259 1380
rect 293 1346 327 1380
rect 361 1346 395 1380
rect 429 1346 463 1380
rect 497 1346 531 1380
rect 565 1346 599 1380
rect 633 1346 667 1380
rect 701 1346 735 1380
rect 769 1346 803 1380
rect 837 1346 871 1380
rect 905 1346 939 1380
rect 973 1346 1007 1380
rect 1041 1346 1075 1380
rect 1109 1346 1143 1380
rect 1177 1346 1211 1380
rect 1245 1346 1279 1380
rect 1313 1346 1347 1380
rect 1381 1346 1415 1380
rect 1449 1346 1483 1380
rect 1517 1346 1551 1380
rect 1585 1346 1619 1380
rect 1653 1346 1687 1380
rect 1721 1346 1755 1380
rect 1789 1346 1823 1380
rect 1857 1346 1891 1380
rect 1925 1346 1959 1380
rect 1993 1346 2027 1380
rect 2061 1346 2095 1380
rect 2129 1346 2163 1380
rect 2197 1346 2231 1380
rect 2265 1346 2299 1380
rect 2333 1346 2367 1380
rect 2401 1346 2435 1380
rect 2469 1346 2503 1380
rect 2537 1346 2571 1380
rect 2605 1346 2639 1380
rect 2673 1346 2707 1380
rect 2741 1346 2775 1380
rect 2809 1346 2843 1380
rect 2877 1346 2911 1380
rect 2945 1346 2979 1380
rect 3013 1346 3047 1380
rect 3081 1346 3115 1380
rect 3149 1346 3196 1380
rect 94 1330 3196 1346
rect 94 1288 194 1330
rect 252 1288 352 1330
rect 410 1288 510 1330
rect 568 1288 668 1330
rect 726 1288 826 1330
rect 884 1288 984 1330
rect 1042 1288 1142 1330
rect 1200 1288 1300 1330
rect 1358 1288 1458 1330
rect 1516 1288 1616 1330
rect 1674 1288 1774 1330
rect 1832 1288 1932 1330
rect 1990 1288 2090 1330
rect 2148 1288 2248 1330
rect 2306 1288 2406 1330
rect 2464 1288 2564 1330
rect 2622 1288 2722 1330
rect 2780 1288 2880 1330
rect 2938 1288 3038 1330
rect 3096 1288 3196 1330
rect 94 -6 194 36
rect 252 -6 352 36
rect 410 -6 510 36
rect 568 -6 668 36
rect 726 -6 826 36
rect 884 -6 984 36
rect 1042 -6 1142 36
rect 1200 -6 1300 36
rect 1358 -6 1458 36
rect 1516 -6 1616 36
rect 1674 -6 1774 36
rect 1832 -6 1932 36
rect 1990 -6 2090 36
rect 2148 -6 2248 36
rect 2306 -6 2406 36
rect 2464 -6 2564 36
rect 2622 -6 2722 36
rect 2780 -6 2880 36
rect 2938 -6 3038 36
rect 3096 -6 3196 36
rect 94 -20 3196 -6
rect 94 -54 123 -20
rect 157 -54 191 -20
rect 225 -54 259 -20
rect 293 -54 327 -20
rect 361 -54 395 -20
rect 429 -54 463 -20
rect 497 -54 531 -20
rect 565 -54 599 -20
rect 633 -54 667 -20
rect 701 -54 735 -20
rect 769 -54 803 -20
rect 837 -54 871 -20
rect 905 -54 939 -20
rect 973 -54 1007 -20
rect 1041 -54 1075 -20
rect 1109 -54 1143 -20
rect 1177 -54 1211 -20
rect 1245 -54 1279 -20
rect 1313 -54 1347 -20
rect 1381 -54 1415 -20
rect 1449 -54 1483 -20
rect 1517 -54 1551 -20
rect 1585 -54 1619 -20
rect 1653 -54 1687 -20
rect 1721 -54 1755 -20
rect 1789 -54 1823 -20
rect 1857 -54 1891 -20
rect 1925 -54 1959 -20
rect 1993 -54 2027 -20
rect 2061 -54 2095 -20
rect 2129 -54 2163 -20
rect 2197 -54 2231 -20
rect 2265 -54 2299 -20
rect 2333 -54 2367 -20
rect 2401 -54 2435 -20
rect 2469 -54 2503 -20
rect 2537 -54 2571 -20
rect 2605 -54 2639 -20
rect 2673 -54 2707 -20
rect 2741 -54 2775 -20
rect 2809 -54 2843 -20
rect 2877 -54 2911 -20
rect 2945 -54 2979 -20
rect 3013 -54 3047 -20
rect 3081 -54 3115 -20
rect 3149 -54 3196 -20
rect 94 -70 3196 -54
<< polycont >>
rect 123 1346 157 1380
rect 191 1346 225 1380
rect 259 1346 293 1380
rect 327 1346 361 1380
rect 395 1346 429 1380
rect 463 1346 497 1380
rect 531 1346 565 1380
rect 599 1346 633 1380
rect 667 1346 701 1380
rect 735 1346 769 1380
rect 803 1346 837 1380
rect 871 1346 905 1380
rect 939 1346 973 1380
rect 1007 1346 1041 1380
rect 1075 1346 1109 1380
rect 1143 1346 1177 1380
rect 1211 1346 1245 1380
rect 1279 1346 1313 1380
rect 1347 1346 1381 1380
rect 1415 1346 1449 1380
rect 1483 1346 1517 1380
rect 1551 1346 1585 1380
rect 1619 1346 1653 1380
rect 1687 1346 1721 1380
rect 1755 1346 1789 1380
rect 1823 1346 1857 1380
rect 1891 1346 1925 1380
rect 1959 1346 1993 1380
rect 2027 1346 2061 1380
rect 2095 1346 2129 1380
rect 2163 1346 2197 1380
rect 2231 1346 2265 1380
rect 2299 1346 2333 1380
rect 2367 1346 2401 1380
rect 2435 1346 2469 1380
rect 2503 1346 2537 1380
rect 2571 1346 2605 1380
rect 2639 1346 2673 1380
rect 2707 1346 2741 1380
rect 2775 1346 2809 1380
rect 2843 1346 2877 1380
rect 2911 1346 2945 1380
rect 2979 1346 3013 1380
rect 3047 1346 3081 1380
rect 3115 1346 3149 1380
rect 123 -54 157 -20
rect 191 -54 225 -20
rect 259 -54 293 -20
rect 327 -54 361 -20
rect 395 -54 429 -20
rect 463 -54 497 -20
rect 531 -54 565 -20
rect 599 -54 633 -20
rect 667 -54 701 -20
rect 735 -54 769 -20
rect 803 -54 837 -20
rect 871 -54 905 -20
rect 939 -54 973 -20
rect 1007 -54 1041 -20
rect 1075 -54 1109 -20
rect 1143 -54 1177 -20
rect 1211 -54 1245 -20
rect 1279 -54 1313 -20
rect 1347 -54 1381 -20
rect 1415 -54 1449 -20
rect 1483 -54 1517 -20
rect 1551 -54 1585 -20
rect 1619 -54 1653 -20
rect 1687 -54 1721 -20
rect 1755 -54 1789 -20
rect 1823 -54 1857 -20
rect 1891 -54 1925 -20
rect 1959 -54 1993 -20
rect 2027 -54 2061 -20
rect 2095 -54 2129 -20
rect 2163 -54 2197 -20
rect 2231 -54 2265 -20
rect 2299 -54 2333 -20
rect 2367 -54 2401 -20
rect 2435 -54 2469 -20
rect 2503 -54 2537 -20
rect 2571 -54 2605 -20
rect 2639 -54 2673 -20
rect 2707 -54 2741 -20
rect 2775 -54 2809 -20
rect 2843 -54 2877 -20
rect 2911 -54 2945 -20
rect 2979 -54 3013 -20
rect 3047 -54 3081 -20
rect 3115 -54 3149 -20
<< locali >>
rect -347 1672 3631 1678
rect -347 1502 152 1672
rect 3178 1502 3631 1672
rect -347 1497 3631 1502
rect -347 1260 -129 1497
rect 94 1380 3196 1394
rect 94 1346 123 1380
rect 177 1346 191 1380
rect 249 1346 259 1380
rect 321 1346 327 1380
rect 393 1346 395 1380
rect 429 1346 431 1380
rect 497 1346 503 1380
rect 565 1346 575 1380
rect 633 1346 647 1380
rect 701 1346 719 1380
rect 769 1346 791 1380
rect 837 1346 863 1380
rect 905 1346 935 1380
rect 973 1346 1007 1380
rect 1041 1346 1075 1380
rect 1113 1346 1143 1380
rect 1185 1346 1211 1380
rect 1257 1346 1279 1380
rect 1329 1346 1347 1380
rect 1401 1346 1415 1380
rect 1473 1346 1483 1380
rect 1545 1346 1551 1380
rect 1617 1346 1619 1380
rect 1653 1346 1655 1380
rect 1721 1346 1727 1380
rect 1789 1346 1799 1380
rect 1857 1346 1871 1380
rect 1925 1346 1943 1380
rect 1993 1346 2015 1380
rect 2061 1346 2087 1380
rect 2129 1346 2159 1380
rect 2197 1346 2231 1380
rect 2265 1346 2299 1380
rect 2337 1346 2367 1380
rect 2409 1346 2435 1380
rect 2481 1346 2503 1380
rect 2553 1346 2571 1380
rect 2625 1346 2639 1380
rect 2697 1346 2707 1380
rect 2769 1346 2775 1380
rect 2841 1346 2843 1380
rect 2877 1346 2879 1380
rect 2945 1346 2951 1380
rect 3013 1346 3023 1380
rect 3081 1346 3095 1380
rect 3149 1346 3196 1380
rect 94 1330 3196 1346
rect -347 657 -323 1260
rect -153 657 -129 1260
rect -347 623 -329 657
rect -151 623 -129 657
rect -347 2 -323 623
rect -153 2 -129 623
rect -347 -184 -129 2
rect 3413 1312 3631 1497
rect 3413 658 3437 1312
rect 3607 658 3631 1312
rect 3413 624 3432 658
rect 3610 624 3631 658
rect 3413 54 3437 624
rect 3607 54 3631 624
rect 94 -20 3196 -6
rect 94 -54 123 -20
rect 177 -54 191 -20
rect 249 -54 259 -20
rect 321 -54 327 -20
rect 393 -54 395 -20
rect 429 -54 431 -20
rect 497 -54 503 -20
rect 565 -54 575 -20
rect 633 -54 647 -20
rect 701 -54 719 -20
rect 769 -54 791 -20
rect 837 -54 863 -20
rect 905 -54 935 -20
rect 973 -54 1007 -20
rect 1041 -54 1075 -20
rect 1113 -54 1143 -20
rect 1185 -54 1211 -20
rect 1257 -54 1279 -20
rect 1329 -54 1347 -20
rect 1401 -54 1415 -20
rect 1473 -54 1483 -20
rect 1545 -54 1551 -20
rect 1617 -54 1619 -20
rect 1653 -54 1655 -20
rect 1721 -54 1727 -20
rect 1789 -54 1799 -20
rect 1857 -54 1871 -20
rect 1925 -54 1943 -20
rect 1993 -54 2015 -20
rect 2061 -54 2087 -20
rect 2129 -54 2159 -20
rect 2197 -54 2231 -20
rect 2265 -54 2299 -20
rect 2337 -54 2367 -20
rect 2409 -54 2435 -20
rect 2481 -54 2503 -20
rect 2553 -54 2571 -20
rect 2625 -54 2639 -20
rect 2697 -54 2707 -20
rect 2769 -54 2775 -20
rect 2841 -54 2843 -20
rect 2877 -54 2879 -20
rect 2945 -54 2951 -20
rect 3013 -54 3023 -20
rect 3081 -54 3095 -20
rect 3149 -54 3196 -20
rect 94 -70 3196 -54
rect 3413 -184 3631 54
rect -347 -190 3631 -184
rect -347 -360 248 -190
rect 3274 -360 3631 -190
rect -347 -365 3631 -360
<< viali >>
rect 143 1346 157 1380
rect 157 1346 177 1380
rect 215 1346 225 1380
rect 225 1346 249 1380
rect 287 1346 293 1380
rect 293 1346 321 1380
rect 359 1346 361 1380
rect 361 1346 393 1380
rect 431 1346 463 1380
rect 463 1346 465 1380
rect 503 1346 531 1380
rect 531 1346 537 1380
rect 575 1346 599 1380
rect 599 1346 609 1380
rect 647 1346 667 1380
rect 667 1346 681 1380
rect 719 1346 735 1380
rect 735 1346 753 1380
rect 791 1346 803 1380
rect 803 1346 825 1380
rect 863 1346 871 1380
rect 871 1346 897 1380
rect 935 1346 939 1380
rect 939 1346 969 1380
rect 1007 1346 1041 1380
rect 1079 1346 1109 1380
rect 1109 1346 1113 1380
rect 1151 1346 1177 1380
rect 1177 1346 1185 1380
rect 1223 1346 1245 1380
rect 1245 1346 1257 1380
rect 1295 1346 1313 1380
rect 1313 1346 1329 1380
rect 1367 1346 1381 1380
rect 1381 1346 1401 1380
rect 1439 1346 1449 1380
rect 1449 1346 1473 1380
rect 1511 1346 1517 1380
rect 1517 1346 1545 1380
rect 1583 1346 1585 1380
rect 1585 1346 1617 1380
rect 1655 1346 1687 1380
rect 1687 1346 1689 1380
rect 1727 1346 1755 1380
rect 1755 1346 1761 1380
rect 1799 1346 1823 1380
rect 1823 1346 1833 1380
rect 1871 1346 1891 1380
rect 1891 1346 1905 1380
rect 1943 1346 1959 1380
rect 1959 1346 1977 1380
rect 2015 1346 2027 1380
rect 2027 1346 2049 1380
rect 2087 1346 2095 1380
rect 2095 1346 2121 1380
rect 2159 1346 2163 1380
rect 2163 1346 2193 1380
rect 2231 1346 2265 1380
rect 2303 1346 2333 1380
rect 2333 1346 2337 1380
rect 2375 1346 2401 1380
rect 2401 1346 2409 1380
rect 2447 1346 2469 1380
rect 2469 1346 2481 1380
rect 2519 1346 2537 1380
rect 2537 1346 2553 1380
rect 2591 1346 2605 1380
rect 2605 1346 2625 1380
rect 2663 1346 2673 1380
rect 2673 1346 2697 1380
rect 2735 1346 2741 1380
rect 2741 1346 2769 1380
rect 2807 1346 2809 1380
rect 2809 1346 2841 1380
rect 2879 1346 2911 1380
rect 2911 1346 2913 1380
rect 2951 1346 2979 1380
rect 2979 1346 2985 1380
rect 3023 1346 3047 1380
rect 3047 1346 3057 1380
rect 3095 1346 3115 1380
rect 3115 1346 3129 1380
rect -329 623 -323 657
rect -323 623 -295 657
rect -257 623 -223 657
rect -185 623 -153 657
rect -153 623 -151 657
rect 3432 624 3437 658
rect 3437 624 3466 658
rect 3504 624 3538 658
rect 3576 624 3607 658
rect 3607 624 3610 658
rect 143 -54 157 -20
rect 157 -54 177 -20
rect 215 -54 225 -20
rect 225 -54 249 -20
rect 287 -54 293 -20
rect 293 -54 321 -20
rect 359 -54 361 -20
rect 361 -54 393 -20
rect 431 -54 463 -20
rect 463 -54 465 -20
rect 503 -54 531 -20
rect 531 -54 537 -20
rect 575 -54 599 -20
rect 599 -54 609 -20
rect 647 -54 667 -20
rect 667 -54 681 -20
rect 719 -54 735 -20
rect 735 -54 753 -20
rect 791 -54 803 -20
rect 803 -54 825 -20
rect 863 -54 871 -20
rect 871 -54 897 -20
rect 935 -54 939 -20
rect 939 -54 969 -20
rect 1007 -54 1041 -20
rect 1079 -54 1109 -20
rect 1109 -54 1113 -20
rect 1151 -54 1177 -20
rect 1177 -54 1185 -20
rect 1223 -54 1245 -20
rect 1245 -54 1257 -20
rect 1295 -54 1313 -20
rect 1313 -54 1329 -20
rect 1367 -54 1381 -20
rect 1381 -54 1401 -20
rect 1439 -54 1449 -20
rect 1449 -54 1473 -20
rect 1511 -54 1517 -20
rect 1517 -54 1545 -20
rect 1583 -54 1585 -20
rect 1585 -54 1617 -20
rect 1655 -54 1687 -20
rect 1687 -54 1689 -20
rect 1727 -54 1755 -20
rect 1755 -54 1761 -20
rect 1799 -54 1823 -20
rect 1823 -54 1833 -20
rect 1871 -54 1891 -20
rect 1891 -54 1905 -20
rect 1943 -54 1959 -20
rect 1959 -54 1977 -20
rect 2015 -54 2027 -20
rect 2027 -54 2049 -20
rect 2087 -54 2095 -20
rect 2095 -54 2121 -20
rect 2159 -54 2163 -20
rect 2163 -54 2193 -20
rect 2231 -54 2265 -20
rect 2303 -54 2333 -20
rect 2333 -54 2337 -20
rect 2375 -54 2401 -20
rect 2401 -54 2409 -20
rect 2447 -54 2469 -20
rect 2469 -54 2481 -20
rect 2519 -54 2537 -20
rect 2537 -54 2553 -20
rect 2591 -54 2605 -20
rect 2605 -54 2625 -20
rect 2663 -54 2673 -20
rect 2673 -54 2697 -20
rect 2735 -54 2741 -20
rect 2741 -54 2769 -20
rect 2807 -54 2809 -20
rect 2809 -54 2841 -20
rect 2879 -54 2911 -20
rect 2911 -54 2913 -20
rect 2951 -54 2979 -20
rect 2979 -54 2985 -20
rect 3023 -54 3047 -20
rect 3047 -54 3057 -20
rect 3095 -54 3115 -20
rect 3115 -54 3129 -20
<< metal1 >>
rect -77 1380 3383 1394
rect -77 1346 143 1380
rect 177 1346 215 1380
rect 249 1346 287 1380
rect 321 1346 359 1380
rect 393 1346 431 1380
rect 465 1346 503 1380
rect 537 1346 575 1380
rect 609 1346 647 1380
rect 681 1346 719 1380
rect 753 1346 791 1380
rect 825 1346 863 1380
rect 897 1346 935 1380
rect 969 1346 1007 1380
rect 1041 1346 1079 1380
rect 1113 1346 1151 1380
rect 1185 1346 1223 1380
rect 1257 1346 1295 1380
rect 1329 1346 1367 1380
rect 1401 1346 1439 1380
rect 1473 1346 1511 1380
rect 1545 1346 1583 1380
rect 1617 1346 1655 1380
rect 1689 1346 1727 1380
rect 1761 1346 1799 1380
rect 1833 1346 1871 1380
rect 1905 1346 1943 1380
rect 1977 1346 2015 1380
rect 2049 1346 2087 1380
rect 2121 1346 2159 1380
rect 2193 1346 2231 1380
rect 2265 1346 2303 1380
rect 2337 1346 2375 1380
rect 2409 1346 2447 1380
rect 2481 1346 2519 1380
rect 2553 1346 2591 1380
rect 2625 1346 2663 1380
rect 2697 1346 2735 1380
rect 2769 1346 2807 1380
rect 2841 1346 2879 1380
rect 2913 1346 2951 1380
rect 2985 1346 3023 1380
rect 3057 1346 3095 1380
rect 3129 1346 3383 1380
rect -77 1330 3383 1346
rect -347 666 -129 698
rect -347 614 -330 666
rect -278 614 -266 666
rect -214 614 -202 666
rect -150 614 -129 666
rect -347 582 -129 614
rect -77 208 -2 1330
rect 349 1187 413 1219
rect 349 1135 355 1187
rect 407 1135 413 1187
rect 349 1103 413 1135
rect 981 1187 1045 1219
rect 981 1135 987 1187
rect 1039 1135 1045 1187
rect 981 1103 1045 1135
rect 1613 1187 1677 1219
rect 1613 1135 1619 1187
rect 1671 1135 1677 1187
rect 1613 1103 1677 1135
rect 2245 1187 2309 1219
rect 2245 1135 2251 1187
rect 2303 1135 2309 1187
rect 2245 1103 2309 1135
rect 2877 1187 2941 1219
rect 2877 1135 2883 1187
rect 2935 1135 2941 1187
rect 2877 1103 2941 1135
rect 191 666 255 698
rect 191 614 197 666
rect 249 614 255 666
rect 191 582 255 614
rect 507 666 571 698
rect 507 614 513 666
rect 565 614 571 666
rect 507 582 571 614
rect 823 666 887 698
rect 823 614 829 666
rect 881 614 887 666
rect 823 582 887 614
rect 1139 666 1203 698
rect 1139 614 1145 666
rect 1197 614 1203 666
rect 1139 582 1203 614
rect 1455 666 1519 698
rect 1455 614 1461 666
rect 1513 614 1519 666
rect 1455 582 1519 614
rect 1771 666 1835 698
rect 1771 614 1777 666
rect 1829 614 1835 666
rect 1771 582 1835 614
rect 2087 666 2151 698
rect 2087 614 2093 666
rect 2145 614 2151 666
rect 2087 582 2151 614
rect 2403 666 2467 698
rect 2403 614 2409 666
rect 2461 614 2467 666
rect 2403 582 2467 614
rect 2719 666 2783 698
rect 2719 614 2725 666
rect 2777 614 2783 666
rect 2719 582 2783 614
rect 3035 666 3099 698
rect 3035 614 3041 666
rect 3093 614 3099 666
rect 3035 582 3099 614
rect 3308 208 3383 1330
rect 3413 667 3631 698
rect 3413 615 3431 667
rect 3483 615 3495 667
rect 3547 615 3559 667
rect 3611 615 3631 667
rect 3413 582 3631 615
rect -77 176 97 208
rect -77 124 39 176
rect 91 124 97 176
rect -77 92 97 124
rect 665 176 729 208
rect 665 124 671 176
rect 723 124 729 176
rect 665 92 729 124
rect 1297 176 1361 208
rect 1297 124 1303 176
rect 1355 124 1361 176
rect 1297 92 1361 124
rect 1929 176 1993 208
rect 1929 124 1935 176
rect 1987 124 1993 176
rect 1929 92 1993 124
rect 2561 176 2625 208
rect 2561 124 2567 176
rect 2619 124 2625 176
rect 2561 92 2625 124
rect 3193 176 3383 208
rect 3193 124 3199 176
rect 3251 124 3383 176
rect 3193 92 3383 124
rect -77 -6 -2 92
rect 3308 -6 3383 92
rect -77 -20 3383 -6
rect -77 -54 143 -20
rect 177 -54 215 -20
rect 249 -54 287 -20
rect 321 -54 359 -20
rect 393 -54 431 -20
rect 465 -54 503 -20
rect 537 -54 575 -20
rect 609 -54 647 -20
rect 681 -54 719 -20
rect 753 -54 791 -20
rect 825 -54 863 -20
rect 897 -54 935 -20
rect 969 -54 1007 -20
rect 1041 -54 1079 -20
rect 1113 -54 1151 -20
rect 1185 -54 1223 -20
rect 1257 -54 1295 -20
rect 1329 -54 1367 -20
rect 1401 -54 1439 -20
rect 1473 -54 1511 -20
rect 1545 -54 1583 -20
rect 1617 -54 1655 -20
rect 1689 -54 1727 -20
rect 1761 -54 1799 -20
rect 1833 -54 1871 -20
rect 1905 -54 1943 -20
rect 1977 -54 2015 -20
rect 2049 -54 2087 -20
rect 2121 -54 2159 -20
rect 2193 -54 2231 -20
rect 2265 -54 2303 -20
rect 2337 -54 2375 -20
rect 2409 -54 2447 -20
rect 2481 -54 2519 -20
rect 2553 -54 2591 -20
rect 2625 -54 2663 -20
rect 2697 -54 2735 -20
rect 2769 -54 2807 -20
rect 2841 -54 2879 -20
rect 2913 -54 2951 -20
rect 2985 -54 3023 -20
rect 3057 -54 3095 -20
rect 3129 -54 3383 -20
rect -77 -70 3383 -54
<< via1 >>
rect -330 657 -278 666
rect -330 623 -329 657
rect -329 623 -295 657
rect -295 623 -278 657
rect -330 614 -278 623
rect -266 657 -214 666
rect -266 623 -257 657
rect -257 623 -223 657
rect -223 623 -214 657
rect -266 614 -214 623
rect -202 657 -150 666
rect -202 623 -185 657
rect -185 623 -151 657
rect -151 623 -150 657
rect -202 614 -150 623
rect 355 1135 407 1187
rect 987 1135 1039 1187
rect 1619 1135 1671 1187
rect 2251 1135 2303 1187
rect 2883 1135 2935 1187
rect 197 614 249 666
rect 513 614 565 666
rect 829 614 881 666
rect 1145 614 1197 666
rect 1461 614 1513 666
rect 1777 614 1829 666
rect 2093 614 2145 666
rect 2409 614 2461 666
rect 2725 614 2777 666
rect 3041 614 3093 666
rect 3431 658 3483 667
rect 3431 624 3432 658
rect 3432 624 3466 658
rect 3466 624 3483 658
rect 3431 615 3483 624
rect 3495 658 3547 667
rect 3495 624 3504 658
rect 3504 624 3538 658
rect 3538 624 3547 658
rect 3495 615 3547 624
rect 3559 658 3611 667
rect 3559 624 3576 658
rect 3576 624 3610 658
rect 3610 624 3611 658
rect 3559 615 3611 624
rect 39 124 91 176
rect 671 124 723 176
rect 1303 124 1355 176
rect 1935 124 1987 176
rect 2567 124 2619 176
rect 3199 124 3251 176
<< metal2 >>
rect -508 1187 3903 1219
rect -508 1135 355 1187
rect 407 1135 987 1187
rect 1039 1135 1619 1187
rect 1671 1135 2251 1187
rect 2303 1135 2883 1187
rect 2935 1135 3903 1187
rect -508 1103 3903 1135
rect -347 667 3631 698
rect -347 666 3431 667
rect -347 614 -330 666
rect -278 614 -266 666
rect -214 614 -202 666
rect -150 614 197 666
rect 249 614 513 666
rect 565 614 829 666
rect 881 614 1145 666
rect 1197 614 1461 666
rect 1513 614 1777 666
rect 1829 614 2093 666
rect 2145 614 2409 666
rect 2461 614 2725 666
rect 2777 614 3041 666
rect 3093 615 3431 666
rect 3483 615 3495 667
rect 3547 615 3559 667
rect 3611 615 3631 667
rect 3093 614 3631 615
rect -347 582 3631 614
rect 36 176 3254 208
rect 36 124 39 176
rect 91 124 671 176
rect 723 124 1303 176
rect 1355 124 1935 176
rect 1987 124 2567 176
rect 2619 124 3199 176
rect 3251 124 3254 176
rect 36 92 3254 124
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_19
timestamp 1640969486
transform 1 0 144 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_18
timestamp 1640969486
transform 1 0 302 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_17
timestamp 1640969486
transform 1 0 460 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_16
timestamp 1640969486
transform 1 0 618 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_15
timestamp 1640969486
transform 1 0 776 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_14
timestamp 1640969486
transform 1 0 934 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_13
timestamp 1640969486
transform 1 0 1092 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_12
timestamp 1640969486
transform 1 0 1250 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_11
timestamp 1640969486
transform 1 0 1408 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_10
timestamp 1640969486
transform 1 0 1566 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_9
timestamp 1640969486
transform 1 0 1724 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_8
timestamp 1640969486
transform 1 0 2040 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_7
timestamp 1640969486
transform 1 0 1882 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_6
timestamp 1640969486
transform 1 0 2356 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_5
timestamp 1640969486
transform 1 0 2198 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_4
timestamp 1640969486
transform 1 0 2672 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_3
timestamp 1640969486
transform 1 0 2514 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_2
timestamp 1640969486
transform 1 0 2988 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_1
timestamp 1640969486
transform 1 0 2830 0 1 662
box -144 -662 144 662
use sky130_fd_pr__pfet_01v8_lvt_EEU9S7  sky130_fd_pr__pfet_01v8_lvt_EEU9S7_0
timestamp 1640969486
transform 1 0 3146 0 1 662
box -144 -662 144 662
<< labels >>
flabel metal2 s -461 1140 -461 1140 0 FreeSans 800 0 0 0 D2
port 1 nsew
flabel metal1 s -53 148 -53 148 0 FreeSans 800 0 0 0 D1
port 2 nsew
flabel metal2 s -100 619 -100 619 0 FreeSans 800 0 0 0 S
port 3 nsew
<< end >>
