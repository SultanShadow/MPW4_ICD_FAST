magic
tech sky130A
magscale 1 2
timestamp 1640969486
<< locali >>
rect 430 9296 504 9334
rect 430 9262 449 9296
rect 483 9262 504 9296
rect 430 9202 504 9262
rect 496 -320 574 -282
rect 496 -354 518 -320
rect 552 -354 574 -320
rect 496 -396 574 -354
rect 16304 -10117 16428 -10040
rect 16304 -10151 16348 -10117
rect 16382 -10151 16428 -10117
rect 16304 -10212 16428 -10151
rect 16268 -19903 16496 -19756
rect 16268 -20081 16332 -19903
rect 16438 -20081 16496 -19903
rect 16268 -20106 16496 -20081
<< viali >>
rect 449 9262 483 9296
rect 518 -354 552 -320
rect 16348 -10151 16382 -10117
rect 16332 -20081 16438 -19903
<< metal1 >>
rect 16366 9344 16582 9474
rect 432 9305 504 9334
rect 432 9253 440 9305
rect 492 9253 504 9305
rect 432 9238 504 9253
rect -14 -176 198 354
rect -14 -228 38 -176
rect 90 -228 102 -176
rect 154 -228 198 -176
rect -14 -248 198 -228
rect 290 144 432 174
rect 290 12 508 144
rect 290 -76 514 12
rect -910 -1034 210 -482
rect 290 -504 432 -76
rect 496 -311 574 -282
rect 496 -363 509 -311
rect 561 -363 574 -311
rect 496 -396 574 -363
rect 74 -9936 272 -9304
rect 74 -10056 606 -9936
rect 16304 -10108 16428 -10040
rect 532 -10216 556 -10130
rect 16304 -10160 16339 -10108
rect 16391 -10160 16428 -10108
rect 16304 -10212 16428 -10160
rect 36 -10436 388 -10336
rect 36 -10552 78 -10436
rect 194 -10552 388 -10436
rect 36 -10642 388 -10552
rect 226 -19826 392 -19276
rect -582 -19888 682 -19826
rect -582 -20004 -561 -19888
rect -381 -20004 682 -19888
rect -582 -20056 682 -20004
rect 16268 -19902 16496 -19756
rect 16268 -20082 16327 -19902
rect 16443 -20082 16496 -19902
rect 16268 -20106 16496 -20082
rect 46 -20294 454 -20246
rect 46 -20474 73 -20294
rect 189 -20474 454 -20294
rect 46 -20498 454 -20474
<< via1 >>
rect 440 9296 492 9305
rect 440 9262 449 9296
rect 449 9262 483 9296
rect 483 9262 492 9296
rect 440 9253 492 9262
rect 38 -228 90 -176
rect 102 -228 154 -176
rect 509 -320 561 -311
rect 509 -354 518 -320
rect 518 -354 552 -320
rect 552 -354 561 -320
rect 509 -363 561 -354
rect 16339 -10117 16391 -10108
rect 16339 -10151 16348 -10117
rect 16348 -10151 16382 -10117
rect 16382 -10151 16391 -10117
rect 16339 -10160 16391 -10151
rect 78 -10552 194 -10436
rect -561 -20004 -381 -19888
rect 16327 -19903 16443 -19902
rect 16327 -20081 16332 -19903
rect 16332 -20081 16438 -19903
rect 16438 -20081 16443 -19903
rect 16327 -20082 16443 -20081
rect 73 -20474 189 -20294
<< metal2 >>
rect 438 9305 494 9308
rect 438 9253 440 9305
rect 492 9253 494 9305
rect 438 9250 494 9253
rect -654 -114 -342 -110
rect -724 -144 224 -114
rect -724 -176 580 -144
rect -724 -228 38 -176
rect 90 -228 102 -176
rect 154 -228 580 -176
rect -724 -248 580 -228
rect -724 -316 224 -248
rect 504 -311 566 -298
rect -654 -19888 -342 -316
rect 504 -363 509 -311
rect 561 -363 566 -311
rect 504 -376 566 -363
rect 16370 -446 16498 440
rect 404 -9654 662 -9382
rect -40 -9664 672 -9654
rect -42 -9862 672 -9664
rect -42 -9908 202 -9862
rect -42 -10436 214 -9908
rect 16292 -10108 17472 -9840
rect 16292 -10156 16339 -10108
rect 16322 -10160 16339 -10156
rect 16391 -10156 17472 -10108
rect 16391 -10160 16408 -10156
rect 16322 -10186 16408 -10160
rect -42 -10444 78 -10436
rect -30 -10552 78 -10444
rect 194 -10450 214 -10436
rect 194 -10552 398 -10450
rect -30 -10688 398 -10552
rect 416 -19582 580 -18916
rect -654 -20004 -561 -19888
rect -381 -20004 -342 -19888
rect -654 -20060 -342 -20004
rect 32 -19770 590 -19582
rect 16270 -19754 16492 -19226
rect 32 -20294 232 -19770
rect 16270 -19902 16496 -19754
rect 16270 -20024 16327 -19902
rect 16276 -20082 16327 -20024
rect 16443 -20082 16496 -19902
rect 16276 -20112 16496 -20082
rect 32 -20474 73 -20294
rect 189 -20474 232 -20294
rect 32 -20498 232 -20474
use pmos20  pmos20_0
timestamp 1640969486
transform 0 1 266 -1 0 9220
box -238 -278 9216 16385
use pmos20  pmos20_1
timestamp 1640969486
transform 0 1 334 -1 0 -342
box -238 -278 9216 16385
use nmos20  nmos20_0
timestamp 1640969486
transform 0 -1 8575 -1 0 -20124
box -308 -8222 9194 8286
use nmos20  nmos20_1
timestamp 1640969486
transform 0 -1 8511 -1 0 -10210
box -308 -8222 9194 8286
<< labels >>
rlabel metal1 s 16536 9384 16536 9384 4 VIN1
port 1 nsew
rlabel metal2 s 17042 -10074 17042 -10074 4 VSS
port 2 nsew
rlabel metal2 s -426 -19954 -426 -19954 4 VINN
port 3 nsew
rlabel metal1 s -146 -846 -146 -846 4 VINP
port 4 nsew
<< end >>
