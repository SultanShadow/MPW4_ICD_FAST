magic
tech sky130A
magscale 1 2
timestamp 1640969486
<< nwell >>
rect 2310 564 8316 579
rect 1289 562 8316 564
rect -917 558 8316 562
rect -1693 549 8316 558
rect -3322 -264 8316 549
rect -3323 -542 8317 -264
<< mvpmos >>
rect 2737 -100 3737 300
rect 3795 -100 4795 300
rect 4853 -100 5853 300
rect 5911 -100 6911 300
rect 6969 -100 7969 300
<< mvpdiff >>
rect 2679 287 2737 300
rect 2679 253 2691 287
rect 2725 253 2737 287
rect 2679 219 2737 253
rect 2679 185 2691 219
rect 2725 185 2737 219
rect 2679 151 2737 185
rect 2679 117 2691 151
rect 2725 117 2737 151
rect 2679 83 2737 117
rect 2679 49 2691 83
rect 2725 49 2737 83
rect 2679 15 2737 49
rect 2679 -19 2691 15
rect 2725 -19 2737 15
rect 2679 -53 2737 -19
rect 2679 -87 2691 -53
rect 2725 -87 2737 -53
rect 2679 -100 2737 -87
rect 3737 287 3795 300
rect 3737 253 3749 287
rect 3783 253 3795 287
rect 3737 219 3795 253
rect 3737 185 3749 219
rect 3783 185 3795 219
rect 3737 151 3795 185
rect 3737 117 3749 151
rect 3783 117 3795 151
rect 3737 83 3795 117
rect 3737 49 3749 83
rect 3783 49 3795 83
rect 3737 15 3795 49
rect 3737 -19 3749 15
rect 3783 -19 3795 15
rect 3737 -53 3795 -19
rect 3737 -87 3749 -53
rect 3783 -87 3795 -53
rect 3737 -100 3795 -87
rect 4795 287 4853 300
rect 4795 253 4807 287
rect 4841 253 4853 287
rect 4795 219 4853 253
rect 4795 185 4807 219
rect 4841 185 4853 219
rect 4795 151 4853 185
rect 4795 117 4807 151
rect 4841 117 4853 151
rect 4795 83 4853 117
rect 4795 49 4807 83
rect 4841 49 4853 83
rect 4795 15 4853 49
rect 4795 -19 4807 15
rect 4841 -19 4853 15
rect 4795 -53 4853 -19
rect 4795 -87 4807 -53
rect 4841 -87 4853 -53
rect 4795 -100 4853 -87
rect 5853 287 5911 300
rect 5853 253 5865 287
rect 5899 253 5911 287
rect 5853 219 5911 253
rect 5853 185 5865 219
rect 5899 185 5911 219
rect 5853 151 5911 185
rect 5853 117 5865 151
rect 5899 117 5911 151
rect 5853 83 5911 117
rect 5853 49 5865 83
rect 5899 49 5911 83
rect 5853 15 5911 49
rect 5853 -19 5865 15
rect 5899 -19 5911 15
rect 5853 -53 5911 -19
rect 5853 -87 5865 -53
rect 5899 -87 5911 -53
rect 5853 -100 5911 -87
rect 6911 287 6969 300
rect 6911 253 6923 287
rect 6957 253 6969 287
rect 6911 219 6969 253
rect 6911 185 6923 219
rect 6957 185 6969 219
rect 6911 151 6969 185
rect 6911 117 6923 151
rect 6957 117 6969 151
rect 6911 83 6969 117
rect 6911 49 6923 83
rect 6957 49 6969 83
rect 6911 15 6969 49
rect 6911 -19 6923 15
rect 6957 -19 6969 15
rect 6911 -53 6969 -19
rect 6911 -87 6923 -53
rect 6957 -87 6969 -53
rect 6911 -100 6969 -87
rect 7969 287 8027 300
rect 7969 253 7981 287
rect 8015 253 8027 287
rect 7969 219 8027 253
rect 7969 185 7981 219
rect 8015 185 8027 219
rect 7969 151 8027 185
rect 7969 117 7981 151
rect 8015 117 8027 151
rect 7969 83 8027 117
rect 7969 49 7981 83
rect 8015 49 8027 83
rect 7969 15 8027 49
rect 7969 -19 7981 15
rect 8015 -19 8027 15
rect 7969 -53 8027 -19
rect 7969 -87 7981 -53
rect 8015 -87 8027 -53
rect 7969 -100 8027 -87
<< mvpdiffc >>
rect 2691 253 2725 287
rect 2691 185 2725 219
rect 2691 117 2725 151
rect 2691 49 2725 83
rect 2691 -19 2725 15
rect 2691 -87 2725 -53
rect 3749 253 3783 287
rect 3749 185 3783 219
rect 3749 117 3783 151
rect 3749 49 3783 83
rect 3749 -19 3783 15
rect 3749 -87 3783 -53
rect 4807 253 4841 287
rect 4807 185 4841 219
rect 4807 117 4841 151
rect 4807 49 4841 83
rect 4807 -19 4841 15
rect 4807 -87 4841 -53
rect 5865 253 5899 287
rect 5865 185 5899 219
rect 5865 117 5899 151
rect 5865 49 5899 83
rect 5865 -19 5899 15
rect 5865 -87 5899 -53
rect 6923 253 6957 287
rect 6923 185 6957 219
rect 6923 117 6957 151
rect 6923 49 6957 83
rect 6923 -19 6957 15
rect 6923 -87 6957 -53
rect 7981 253 8015 287
rect 7981 185 8015 219
rect 7981 117 8015 151
rect 7981 49 8015 83
rect 7981 -19 8015 15
rect 7981 -87 8015 -53
<< poly >>
rect 2333 497 2757 509
rect 2333 482 7967 497
rect -2894 477 7967 482
rect -2894 462 2786 477
rect -2894 428 -2844 462
rect -2810 428 -2776 462
rect -2742 428 -2708 462
rect -2674 428 -2640 462
rect -2606 428 -2572 462
rect -2538 428 -2504 462
rect -2470 428 -2436 462
rect -2402 428 -2368 462
rect -2334 428 -2300 462
rect -2266 428 -2232 462
rect -2198 428 -2164 462
rect -2130 428 -2096 462
rect -2062 428 -2028 462
rect -1994 428 -1960 462
rect -1926 428 -1892 462
rect -1858 428 -1824 462
rect -1790 428 -1756 462
rect -1722 428 -1688 462
rect -1654 428 -1620 462
rect -1586 428 -1552 462
rect -1518 428 -1484 462
rect -1450 428 -1416 462
rect -1382 428 -1348 462
rect -1314 428 -1280 462
rect -1246 428 -1212 462
rect -1178 428 -1144 462
rect -1110 428 -1076 462
rect -1042 428 -1008 462
rect -974 428 -940 462
rect -906 428 -872 462
rect -838 428 -804 462
rect -770 428 -736 462
rect -702 428 -668 462
rect -634 428 -600 462
rect -566 428 -532 462
rect -498 428 -464 462
rect -430 428 -396 462
rect -362 428 -328 462
rect -294 428 -260 462
rect -226 428 -192 462
rect -158 428 -124 462
rect -90 428 -56 462
rect -22 428 12 462
rect 46 428 80 462
rect 114 428 148 462
rect 182 428 216 462
rect 250 428 284 462
rect 318 428 352 462
rect 386 428 420 462
rect 454 428 488 462
rect 522 428 556 462
rect 590 428 624 462
rect 658 428 692 462
rect 726 428 760 462
rect 794 428 828 462
rect 862 428 896 462
rect 930 428 964 462
rect 998 428 1032 462
rect 1066 428 1100 462
rect 1134 428 1168 462
rect 1202 428 1236 462
rect 1270 428 1304 462
rect 1338 428 1372 462
rect 1406 428 1440 462
rect 1474 428 1508 462
rect 1542 428 1576 462
rect 1610 428 1644 462
rect 1678 428 1712 462
rect 1746 428 1780 462
rect 1814 428 1848 462
rect 1882 428 1916 462
rect 1950 428 1984 462
rect 2018 428 2052 462
rect 2086 428 2120 462
rect 2154 428 2188 462
rect 2222 428 2256 462
rect 2290 443 2786 462
rect 2820 443 2854 477
rect 2888 443 2922 477
rect 2956 443 2990 477
rect 3024 443 3058 477
rect 3092 443 3126 477
rect 3160 443 3194 477
rect 3228 443 3262 477
rect 3296 443 3330 477
rect 3364 443 3398 477
rect 3432 443 3466 477
rect 3500 443 3534 477
rect 3568 443 3602 477
rect 3636 443 3670 477
rect 3704 443 3738 477
rect 3772 443 3806 477
rect 3840 443 3874 477
rect 3908 443 3942 477
rect 3976 443 4010 477
rect 4044 443 4078 477
rect 4112 443 4146 477
rect 4180 443 4214 477
rect 4248 443 4282 477
rect 4316 443 4350 477
rect 4384 443 4418 477
rect 4452 443 4486 477
rect 4520 443 4554 477
rect 4588 443 4622 477
rect 4656 443 4690 477
rect 4724 443 4758 477
rect 4792 443 4826 477
rect 4860 443 4894 477
rect 4928 443 4962 477
rect 4996 443 5030 477
rect 5064 443 5098 477
rect 5132 443 5166 477
rect 5200 443 5234 477
rect 5268 443 5302 477
rect 5336 443 5370 477
rect 5404 443 5438 477
rect 5472 443 5506 477
rect 5540 443 5574 477
rect 5608 443 5642 477
rect 5676 443 5710 477
rect 5744 443 5778 477
rect 5812 443 5846 477
rect 5880 443 5914 477
rect 5948 443 5982 477
rect 6016 443 6050 477
rect 6084 443 6118 477
rect 6152 443 6186 477
rect 6220 443 6254 477
rect 6288 443 6322 477
rect 6356 443 6390 477
rect 6424 443 6458 477
rect 6492 443 6526 477
rect 6560 443 6594 477
rect 6628 443 6662 477
rect 6696 443 6730 477
rect 6764 443 6798 477
rect 6832 443 6866 477
rect 6900 443 6934 477
rect 6968 443 7002 477
rect 7036 443 7070 477
rect 7104 443 7138 477
rect 7172 443 7206 477
rect 7240 443 7274 477
rect 7308 443 7342 477
rect 7376 443 7410 477
rect 7444 443 7478 477
rect 7512 443 7546 477
rect 7580 443 7614 477
rect 7648 443 7682 477
rect 7716 443 7750 477
rect 7784 443 7818 477
rect 7852 443 7886 477
rect 7920 443 7967 477
rect 2290 428 7967 443
rect -2894 422 7967 428
rect -2894 419 7968 422
rect -2894 404 3736 419
rect -2894 311 -1894 404
rect -1836 311 -836 404
rect -778 311 222 404
rect 280 311 1280 404
rect 1338 403 3736 404
rect 1338 311 2338 403
rect 2736 326 3736 403
rect 3794 326 4794 419
rect 4852 326 5852 419
rect 5910 326 6910 419
rect 6968 326 7968 419
rect 2737 300 3737 326
rect 3795 300 4795 326
rect 4853 300 5853 326
rect 5911 300 6911 326
rect 6969 300 7969 326
rect 2737 -126 3737 -100
rect 3795 -126 4795 -100
rect 4853 -126 5853 -100
rect 5911 -126 6911 -100
rect 6969 -126 7969 -100
<< polycont >>
rect -2844 428 -2810 462
rect -2776 428 -2742 462
rect -2708 428 -2674 462
rect -2640 428 -2606 462
rect -2572 428 -2538 462
rect -2504 428 -2470 462
rect -2436 428 -2402 462
rect -2368 428 -2334 462
rect -2300 428 -2266 462
rect -2232 428 -2198 462
rect -2164 428 -2130 462
rect -2096 428 -2062 462
rect -2028 428 -1994 462
rect -1960 428 -1926 462
rect -1892 428 -1858 462
rect -1824 428 -1790 462
rect -1756 428 -1722 462
rect -1688 428 -1654 462
rect -1620 428 -1586 462
rect -1552 428 -1518 462
rect -1484 428 -1450 462
rect -1416 428 -1382 462
rect -1348 428 -1314 462
rect -1280 428 -1246 462
rect -1212 428 -1178 462
rect -1144 428 -1110 462
rect -1076 428 -1042 462
rect -1008 428 -974 462
rect -940 428 -906 462
rect -872 428 -838 462
rect -804 428 -770 462
rect -736 428 -702 462
rect -668 428 -634 462
rect -600 428 -566 462
rect -532 428 -498 462
rect -464 428 -430 462
rect -396 428 -362 462
rect -328 428 -294 462
rect -260 428 -226 462
rect -192 428 -158 462
rect -124 428 -90 462
rect -56 428 -22 462
rect 12 428 46 462
rect 80 428 114 462
rect 148 428 182 462
rect 216 428 250 462
rect 284 428 318 462
rect 352 428 386 462
rect 420 428 454 462
rect 488 428 522 462
rect 556 428 590 462
rect 624 428 658 462
rect 692 428 726 462
rect 760 428 794 462
rect 828 428 862 462
rect 896 428 930 462
rect 964 428 998 462
rect 1032 428 1066 462
rect 1100 428 1134 462
rect 1168 428 1202 462
rect 1236 428 1270 462
rect 1304 428 1338 462
rect 1372 428 1406 462
rect 1440 428 1474 462
rect 1508 428 1542 462
rect 1576 428 1610 462
rect 1644 428 1678 462
rect 1712 428 1746 462
rect 1780 428 1814 462
rect 1848 428 1882 462
rect 1916 428 1950 462
rect 1984 428 2018 462
rect 2052 428 2086 462
rect 2120 428 2154 462
rect 2188 428 2222 462
rect 2256 428 2290 462
rect 2786 443 2820 477
rect 2854 443 2888 477
rect 2922 443 2956 477
rect 2990 443 3024 477
rect 3058 443 3092 477
rect 3126 443 3160 477
rect 3194 443 3228 477
rect 3262 443 3296 477
rect 3330 443 3364 477
rect 3398 443 3432 477
rect 3466 443 3500 477
rect 3534 443 3568 477
rect 3602 443 3636 477
rect 3670 443 3704 477
rect 3738 443 3772 477
rect 3806 443 3840 477
rect 3874 443 3908 477
rect 3942 443 3976 477
rect 4010 443 4044 477
rect 4078 443 4112 477
rect 4146 443 4180 477
rect 4214 443 4248 477
rect 4282 443 4316 477
rect 4350 443 4384 477
rect 4418 443 4452 477
rect 4486 443 4520 477
rect 4554 443 4588 477
rect 4622 443 4656 477
rect 4690 443 4724 477
rect 4758 443 4792 477
rect 4826 443 4860 477
rect 4894 443 4928 477
rect 4962 443 4996 477
rect 5030 443 5064 477
rect 5098 443 5132 477
rect 5166 443 5200 477
rect 5234 443 5268 477
rect 5302 443 5336 477
rect 5370 443 5404 477
rect 5438 443 5472 477
rect 5506 443 5540 477
rect 5574 443 5608 477
rect 5642 443 5676 477
rect 5710 443 5744 477
rect 5778 443 5812 477
rect 5846 443 5880 477
rect 5914 443 5948 477
rect 5982 443 6016 477
rect 6050 443 6084 477
rect 6118 443 6152 477
rect 6186 443 6220 477
rect 6254 443 6288 477
rect 6322 443 6356 477
rect 6390 443 6424 477
rect 6458 443 6492 477
rect 6526 443 6560 477
rect 6594 443 6628 477
rect 6662 443 6696 477
rect 6730 443 6764 477
rect 6798 443 6832 477
rect 6866 443 6900 477
rect 6934 443 6968 477
rect 7002 443 7036 477
rect 7070 443 7104 477
rect 7138 443 7172 477
rect 7206 443 7240 477
rect 7274 443 7308 477
rect 7342 443 7376 477
rect 7410 443 7444 477
rect 7478 443 7512 477
rect 7546 443 7580 477
rect 7614 443 7648 477
rect 7682 443 7716 477
rect 7750 443 7784 477
rect 7818 443 7852 477
rect 7886 443 7920 477
<< locali >>
rect 2333 497 2757 509
rect 2333 482 7967 497
rect -2894 477 7967 482
rect -2894 462 2779 477
rect -2894 428 -2851 462
rect -2810 428 -2779 462
rect -2742 428 -2708 462
rect -2673 428 -2640 462
rect -2601 428 -2572 462
rect -2529 428 -2504 462
rect -2457 428 -2436 462
rect -2385 428 -2368 462
rect -2313 428 -2300 462
rect -2241 428 -2232 462
rect -2169 428 -2164 462
rect -2097 428 -2096 462
rect -2062 428 -2059 462
rect -1994 428 -1987 462
rect -1926 428 -1915 462
rect -1858 428 -1843 462
rect -1790 428 -1771 462
rect -1722 428 -1699 462
rect -1654 428 -1627 462
rect -1586 428 -1555 462
rect -1518 428 -1484 462
rect -1449 428 -1416 462
rect -1377 428 -1348 462
rect -1305 428 -1280 462
rect -1233 428 -1212 462
rect -1161 428 -1144 462
rect -1089 428 -1076 462
rect -1017 428 -1008 462
rect -945 428 -940 462
rect -873 428 -872 462
rect -838 428 -835 462
rect -770 428 -763 462
rect -702 428 -691 462
rect -634 428 -619 462
rect -566 428 -547 462
rect -498 428 -475 462
rect -430 428 -403 462
rect -362 428 -331 462
rect -294 428 -260 462
rect -225 428 -192 462
rect -153 428 -124 462
rect -81 428 -56 462
rect -9 428 12 462
rect 63 428 80 462
rect 135 428 148 462
rect 207 428 216 462
rect 279 428 284 462
rect 351 428 352 462
rect 386 428 389 462
rect 454 428 461 462
rect 522 428 533 462
rect 590 428 605 462
rect 658 428 677 462
rect 726 428 749 462
rect 794 428 821 462
rect 862 428 893 462
rect 930 428 964 462
rect 999 428 1032 462
rect 1071 428 1100 462
rect 1143 428 1168 462
rect 1215 428 1236 462
rect 1287 428 1304 462
rect 1359 428 1372 462
rect 1431 428 1440 462
rect 1503 428 1508 462
rect 1575 428 1576 462
rect 1610 428 1613 462
rect 1678 428 1685 462
rect 1746 428 1757 462
rect 1814 428 1829 462
rect 1882 428 1901 462
rect 1950 428 1973 462
rect 2018 428 2045 462
rect 2086 428 2117 462
rect 2154 428 2188 462
rect 2223 428 2256 462
rect 2295 443 2779 462
rect 2820 443 2851 477
rect 2888 443 2922 477
rect 2957 443 2990 477
rect 3029 443 3058 477
rect 3101 443 3126 477
rect 3173 443 3194 477
rect 3245 443 3262 477
rect 3317 443 3330 477
rect 3389 443 3398 477
rect 3461 443 3466 477
rect 3533 443 3534 477
rect 3568 443 3571 477
rect 3636 443 3643 477
rect 3704 443 3715 477
rect 3772 443 3787 477
rect 3840 443 3859 477
rect 3908 443 3931 477
rect 3976 443 4003 477
rect 4044 443 4075 477
rect 4112 443 4146 477
rect 4181 443 4214 477
rect 4253 443 4282 477
rect 4325 443 4350 477
rect 4397 443 4418 477
rect 4469 443 4486 477
rect 4541 443 4554 477
rect 4613 443 4622 477
rect 4685 443 4690 477
rect 4757 443 4758 477
rect 4792 443 4795 477
rect 4860 443 4867 477
rect 4928 443 4939 477
rect 4996 443 5011 477
rect 5064 443 5083 477
rect 5132 443 5155 477
rect 5200 443 5227 477
rect 5268 443 5299 477
rect 5336 443 5370 477
rect 5405 443 5438 477
rect 5477 443 5506 477
rect 5549 443 5574 477
rect 5621 443 5642 477
rect 5693 443 5710 477
rect 5765 443 5778 477
rect 5837 443 5846 477
rect 5909 443 5914 477
rect 5981 443 5982 477
rect 6016 443 6019 477
rect 6084 443 6091 477
rect 6152 443 6163 477
rect 6220 443 6235 477
rect 6288 443 6307 477
rect 6356 443 6379 477
rect 6424 443 6451 477
rect 6492 443 6523 477
rect 6560 443 6594 477
rect 6629 443 6662 477
rect 6701 443 6730 477
rect 6773 443 6798 477
rect 6845 443 6866 477
rect 6917 443 6934 477
rect 6989 443 7002 477
rect 7061 443 7070 477
rect 7133 443 7138 477
rect 7205 443 7206 477
rect 7240 443 7243 477
rect 7308 443 7315 477
rect 7376 443 7387 477
rect 7444 443 7459 477
rect 7512 443 7531 477
rect 7580 443 7603 477
rect 7648 443 7675 477
rect 7716 443 7747 477
rect 7784 443 7818 477
rect 7853 443 7886 477
rect 7925 443 7967 477
rect 2295 428 7967 443
rect -2894 417 7967 428
rect -2894 403 2757 417
rect -2894 402 2337 403
rect 2691 287 2725 304
rect 2691 219 2725 227
rect 2691 151 2725 155
rect 2691 45 2725 49
rect 2691 -27 2725 -19
rect -2939 -173 -2905 -118
rect -823 -173 -789 -118
rect 1293 -173 1327 -118
rect 2691 -158 2725 -87
rect 3749 287 3783 304
rect 3749 219 3783 227
rect 3749 151 3783 155
rect 3749 45 3783 49
rect 3749 -27 3783 -19
rect 3749 -104 3783 -87
rect 4807 287 4841 304
rect 4807 219 4841 227
rect 4807 151 4841 155
rect 4807 45 4841 49
rect 4807 -27 4841 -19
rect 4807 -158 4841 -87
rect 5865 287 5899 304
rect 5865 219 5899 227
rect 5865 151 5899 155
rect 5865 45 5899 49
rect 5865 -27 5899 -19
rect 5865 -104 5899 -87
rect 6923 287 6957 304
rect 6923 219 6957 227
rect 6923 151 6957 155
rect 6923 45 6957 49
rect 6923 -27 6957 -19
rect 6923 -158 6957 -87
rect 7981 287 8015 304
rect 7981 219 8015 227
rect 7981 151 8015 155
rect 7981 45 8015 49
rect 7981 -27 8015 -19
rect 7981 -104 8015 -87
rect 2691 -159 6958 -158
rect -2939 -217 1328 -173
rect 2688 -202 6958 -159
rect 1127 -298 1327 -217
rect 2688 -297 2976 -202
rect 3750 -297 4005 -202
rect 2252 -298 4006 -297
rect 1127 -445 4007 -298
rect 1127 -446 2981 -445
<< viali >>
rect -2851 428 -2844 462
rect -2844 428 -2817 462
rect -2779 428 -2776 462
rect -2776 428 -2745 462
rect -2707 428 -2674 462
rect -2674 428 -2673 462
rect -2635 428 -2606 462
rect -2606 428 -2601 462
rect -2563 428 -2538 462
rect -2538 428 -2529 462
rect -2491 428 -2470 462
rect -2470 428 -2457 462
rect -2419 428 -2402 462
rect -2402 428 -2385 462
rect -2347 428 -2334 462
rect -2334 428 -2313 462
rect -2275 428 -2266 462
rect -2266 428 -2241 462
rect -2203 428 -2198 462
rect -2198 428 -2169 462
rect -2131 428 -2130 462
rect -2130 428 -2097 462
rect -2059 428 -2028 462
rect -2028 428 -2025 462
rect -1987 428 -1960 462
rect -1960 428 -1953 462
rect -1915 428 -1892 462
rect -1892 428 -1881 462
rect -1843 428 -1824 462
rect -1824 428 -1809 462
rect -1771 428 -1756 462
rect -1756 428 -1737 462
rect -1699 428 -1688 462
rect -1688 428 -1665 462
rect -1627 428 -1620 462
rect -1620 428 -1593 462
rect -1555 428 -1552 462
rect -1552 428 -1521 462
rect -1483 428 -1450 462
rect -1450 428 -1449 462
rect -1411 428 -1382 462
rect -1382 428 -1377 462
rect -1339 428 -1314 462
rect -1314 428 -1305 462
rect -1267 428 -1246 462
rect -1246 428 -1233 462
rect -1195 428 -1178 462
rect -1178 428 -1161 462
rect -1123 428 -1110 462
rect -1110 428 -1089 462
rect -1051 428 -1042 462
rect -1042 428 -1017 462
rect -979 428 -974 462
rect -974 428 -945 462
rect -907 428 -906 462
rect -906 428 -873 462
rect -835 428 -804 462
rect -804 428 -801 462
rect -763 428 -736 462
rect -736 428 -729 462
rect -691 428 -668 462
rect -668 428 -657 462
rect -619 428 -600 462
rect -600 428 -585 462
rect -547 428 -532 462
rect -532 428 -513 462
rect -475 428 -464 462
rect -464 428 -441 462
rect -403 428 -396 462
rect -396 428 -369 462
rect -331 428 -328 462
rect -328 428 -297 462
rect -259 428 -226 462
rect -226 428 -225 462
rect -187 428 -158 462
rect -158 428 -153 462
rect -115 428 -90 462
rect -90 428 -81 462
rect -43 428 -22 462
rect -22 428 -9 462
rect 29 428 46 462
rect 46 428 63 462
rect 101 428 114 462
rect 114 428 135 462
rect 173 428 182 462
rect 182 428 207 462
rect 245 428 250 462
rect 250 428 279 462
rect 317 428 318 462
rect 318 428 351 462
rect 389 428 420 462
rect 420 428 423 462
rect 461 428 488 462
rect 488 428 495 462
rect 533 428 556 462
rect 556 428 567 462
rect 605 428 624 462
rect 624 428 639 462
rect 677 428 692 462
rect 692 428 711 462
rect 749 428 760 462
rect 760 428 783 462
rect 821 428 828 462
rect 828 428 855 462
rect 893 428 896 462
rect 896 428 927 462
rect 965 428 998 462
rect 998 428 999 462
rect 1037 428 1066 462
rect 1066 428 1071 462
rect 1109 428 1134 462
rect 1134 428 1143 462
rect 1181 428 1202 462
rect 1202 428 1215 462
rect 1253 428 1270 462
rect 1270 428 1287 462
rect 1325 428 1338 462
rect 1338 428 1359 462
rect 1397 428 1406 462
rect 1406 428 1431 462
rect 1469 428 1474 462
rect 1474 428 1503 462
rect 1541 428 1542 462
rect 1542 428 1575 462
rect 1613 428 1644 462
rect 1644 428 1647 462
rect 1685 428 1712 462
rect 1712 428 1719 462
rect 1757 428 1780 462
rect 1780 428 1791 462
rect 1829 428 1848 462
rect 1848 428 1863 462
rect 1901 428 1916 462
rect 1916 428 1935 462
rect 1973 428 1984 462
rect 1984 428 2007 462
rect 2045 428 2052 462
rect 2052 428 2079 462
rect 2117 428 2120 462
rect 2120 428 2151 462
rect 2189 428 2222 462
rect 2222 428 2223 462
rect 2261 428 2290 462
rect 2290 428 2295 462
rect 2779 443 2786 477
rect 2786 443 2813 477
rect 2851 443 2854 477
rect 2854 443 2885 477
rect 2923 443 2956 477
rect 2956 443 2957 477
rect 2995 443 3024 477
rect 3024 443 3029 477
rect 3067 443 3092 477
rect 3092 443 3101 477
rect 3139 443 3160 477
rect 3160 443 3173 477
rect 3211 443 3228 477
rect 3228 443 3245 477
rect 3283 443 3296 477
rect 3296 443 3317 477
rect 3355 443 3364 477
rect 3364 443 3389 477
rect 3427 443 3432 477
rect 3432 443 3461 477
rect 3499 443 3500 477
rect 3500 443 3533 477
rect 3571 443 3602 477
rect 3602 443 3605 477
rect 3643 443 3670 477
rect 3670 443 3677 477
rect 3715 443 3738 477
rect 3738 443 3749 477
rect 3787 443 3806 477
rect 3806 443 3821 477
rect 3859 443 3874 477
rect 3874 443 3893 477
rect 3931 443 3942 477
rect 3942 443 3965 477
rect 4003 443 4010 477
rect 4010 443 4037 477
rect 4075 443 4078 477
rect 4078 443 4109 477
rect 4147 443 4180 477
rect 4180 443 4181 477
rect 4219 443 4248 477
rect 4248 443 4253 477
rect 4291 443 4316 477
rect 4316 443 4325 477
rect 4363 443 4384 477
rect 4384 443 4397 477
rect 4435 443 4452 477
rect 4452 443 4469 477
rect 4507 443 4520 477
rect 4520 443 4541 477
rect 4579 443 4588 477
rect 4588 443 4613 477
rect 4651 443 4656 477
rect 4656 443 4685 477
rect 4723 443 4724 477
rect 4724 443 4757 477
rect 4795 443 4826 477
rect 4826 443 4829 477
rect 4867 443 4894 477
rect 4894 443 4901 477
rect 4939 443 4962 477
rect 4962 443 4973 477
rect 5011 443 5030 477
rect 5030 443 5045 477
rect 5083 443 5098 477
rect 5098 443 5117 477
rect 5155 443 5166 477
rect 5166 443 5189 477
rect 5227 443 5234 477
rect 5234 443 5261 477
rect 5299 443 5302 477
rect 5302 443 5333 477
rect 5371 443 5404 477
rect 5404 443 5405 477
rect 5443 443 5472 477
rect 5472 443 5477 477
rect 5515 443 5540 477
rect 5540 443 5549 477
rect 5587 443 5608 477
rect 5608 443 5621 477
rect 5659 443 5676 477
rect 5676 443 5693 477
rect 5731 443 5744 477
rect 5744 443 5765 477
rect 5803 443 5812 477
rect 5812 443 5837 477
rect 5875 443 5880 477
rect 5880 443 5909 477
rect 5947 443 5948 477
rect 5948 443 5981 477
rect 6019 443 6050 477
rect 6050 443 6053 477
rect 6091 443 6118 477
rect 6118 443 6125 477
rect 6163 443 6186 477
rect 6186 443 6197 477
rect 6235 443 6254 477
rect 6254 443 6269 477
rect 6307 443 6322 477
rect 6322 443 6341 477
rect 6379 443 6390 477
rect 6390 443 6413 477
rect 6451 443 6458 477
rect 6458 443 6485 477
rect 6523 443 6526 477
rect 6526 443 6557 477
rect 6595 443 6628 477
rect 6628 443 6629 477
rect 6667 443 6696 477
rect 6696 443 6701 477
rect 6739 443 6764 477
rect 6764 443 6773 477
rect 6811 443 6832 477
rect 6832 443 6845 477
rect 6883 443 6900 477
rect 6900 443 6917 477
rect 6955 443 6968 477
rect 6968 443 6989 477
rect 7027 443 7036 477
rect 7036 443 7061 477
rect 7099 443 7104 477
rect 7104 443 7133 477
rect 7171 443 7172 477
rect 7172 443 7205 477
rect 7243 443 7274 477
rect 7274 443 7277 477
rect 7315 443 7342 477
rect 7342 443 7349 477
rect 7387 443 7410 477
rect 7410 443 7421 477
rect 7459 443 7478 477
rect 7478 443 7493 477
rect 7531 443 7546 477
rect 7546 443 7565 477
rect 7603 443 7614 477
rect 7614 443 7637 477
rect 7675 443 7682 477
rect 7682 443 7709 477
rect 7747 443 7750 477
rect 7750 443 7781 477
rect 7819 443 7852 477
rect 7852 443 7853 477
rect 7891 443 7920 477
rect 7920 443 7925 477
rect 2691 253 2725 261
rect 2691 227 2725 253
rect 2691 185 2725 189
rect 2691 155 2725 185
rect 2691 83 2725 117
rect 2691 15 2725 45
rect 2691 11 2725 15
rect 2691 -53 2725 -27
rect 2691 -61 2725 -53
rect 3749 253 3783 261
rect 3749 227 3783 253
rect 3749 185 3783 189
rect 3749 155 3783 185
rect 3749 83 3783 117
rect 3749 15 3783 45
rect 3749 11 3783 15
rect 3749 -53 3783 -27
rect 3749 -61 3783 -53
rect 4807 253 4841 261
rect 4807 227 4841 253
rect 4807 185 4841 189
rect 4807 155 4841 185
rect 4807 83 4841 117
rect 4807 15 4841 45
rect 4807 11 4841 15
rect 4807 -53 4841 -27
rect 4807 -61 4841 -53
rect 5865 253 5899 261
rect 5865 227 5899 253
rect 5865 185 5899 189
rect 5865 155 5899 185
rect 5865 83 5899 117
rect 5865 15 5899 45
rect 5865 11 5899 15
rect 5865 -53 5899 -27
rect 5865 -61 5899 -53
rect 6923 253 6957 261
rect 6923 227 6957 253
rect 6923 185 6957 189
rect 6923 155 6957 185
rect 6923 83 6957 117
rect 6923 15 6957 45
rect 6923 11 6957 15
rect 6923 -53 6957 -27
rect 6923 -61 6957 -53
rect 7981 253 8015 261
rect 7981 227 8015 253
rect 7981 185 8015 189
rect 7981 155 8015 185
rect 7981 83 8015 117
rect 7981 15 8015 45
rect 7981 11 8015 15
rect 7981 -53 8015 -27
rect 7981 -61 8015 -53
<< metal1 >>
rect 2333 497 2757 509
rect 2333 482 7967 497
rect -2894 477 7967 482
rect -2894 462 2779 477
rect -2894 428 -2851 462
rect -2817 428 -2779 462
rect -2745 428 -2707 462
rect -2673 428 -2635 462
rect -2601 428 -2563 462
rect -2529 428 -2491 462
rect -2457 428 -2419 462
rect -2385 428 -2347 462
rect -2313 428 -2275 462
rect -2241 428 -2203 462
rect -2169 428 -2131 462
rect -2097 428 -2059 462
rect -2025 428 -1987 462
rect -1953 428 -1915 462
rect -1881 428 -1843 462
rect -1809 428 -1771 462
rect -1737 428 -1699 462
rect -1665 428 -1627 462
rect -1593 428 -1555 462
rect -1521 428 -1483 462
rect -1449 428 -1411 462
rect -1377 428 -1339 462
rect -1305 428 -1267 462
rect -1233 428 -1195 462
rect -1161 428 -1123 462
rect -1089 428 -1051 462
rect -1017 428 -979 462
rect -945 428 -907 462
rect -873 428 -835 462
rect -801 428 -763 462
rect -729 428 -691 462
rect -657 428 -619 462
rect -585 428 -547 462
rect -513 428 -475 462
rect -441 428 -403 462
rect -369 428 -331 462
rect -297 428 -259 462
rect -225 428 -187 462
rect -153 428 -115 462
rect -81 428 -43 462
rect -9 428 29 462
rect 63 428 101 462
rect 135 428 173 462
rect 207 428 245 462
rect 279 428 317 462
rect 351 428 389 462
rect 423 428 461 462
rect 495 428 533 462
rect 567 428 605 462
rect 639 428 677 462
rect 711 428 749 462
rect 783 428 821 462
rect 855 428 893 462
rect 927 428 965 462
rect 999 428 1037 462
rect 1071 428 1109 462
rect 1143 428 1181 462
rect 1215 428 1253 462
rect 1287 428 1325 462
rect 1359 428 1397 462
rect 1431 428 1469 462
rect 1503 428 1541 462
rect 1575 428 1613 462
rect 1647 428 1685 462
rect 1719 428 1757 462
rect 1791 428 1829 462
rect 1863 428 1901 462
rect 1935 428 1973 462
rect 2007 428 2045 462
rect 2079 428 2117 462
rect 2151 428 2189 462
rect 2223 428 2261 462
rect 2295 443 2779 462
rect 2813 443 2851 477
rect 2885 443 2923 477
rect 2957 443 2995 477
rect 3029 443 3067 477
rect 3101 443 3139 477
rect 3173 443 3211 477
rect 3245 443 3283 477
rect 3317 443 3355 477
rect 3389 443 3427 477
rect 3461 443 3499 477
rect 3533 443 3571 477
rect 3605 443 3643 477
rect 3677 443 3715 477
rect 3749 443 3787 477
rect 3821 443 3859 477
rect 3893 443 3931 477
rect 3965 443 4003 477
rect 4037 443 4075 477
rect 4109 443 4147 477
rect 4181 443 4219 477
rect 4253 443 4291 477
rect 4325 443 4363 477
rect 4397 443 4435 477
rect 4469 443 4507 477
rect 4541 443 4579 477
rect 4613 443 4651 477
rect 4685 443 4723 477
rect 4757 443 4795 477
rect 4829 443 4867 477
rect 4901 443 4939 477
rect 4973 443 5011 477
rect 5045 443 5083 477
rect 5117 443 5155 477
rect 5189 443 5227 477
rect 5261 443 5299 477
rect 5333 443 5371 477
rect 5405 443 5443 477
rect 5477 443 5515 477
rect 5549 443 5587 477
rect 5621 443 5659 477
rect 5693 443 5731 477
rect 5765 443 5803 477
rect 5837 443 5875 477
rect 5909 443 5947 477
rect 5981 443 6019 477
rect 6053 443 6091 477
rect 6125 443 6163 477
rect 6197 443 6235 477
rect 6269 443 6307 477
rect 6341 443 6379 477
rect 6413 443 6451 477
rect 6485 443 6523 477
rect 6557 443 6595 477
rect 6629 443 6667 477
rect 6701 443 6739 477
rect 6773 443 6811 477
rect 6845 443 6883 477
rect 6917 443 6955 477
rect 6989 443 7027 477
rect 7061 443 7099 477
rect 7133 443 7171 477
rect 7205 443 7243 477
rect 7277 443 7315 477
rect 7349 443 7387 477
rect 7421 443 7459 477
rect 7493 443 7531 477
rect 7565 443 7603 477
rect 7637 443 7675 477
rect 7709 443 7747 477
rect 7781 443 7819 477
rect 7853 443 7891 477
rect 7925 443 7967 477
rect 2295 428 7967 443
rect -2894 417 7967 428
rect -2894 403 2757 417
rect -2894 402 2337 403
rect 2685 261 2731 300
rect 2685 227 2691 261
rect 2725 227 2731 261
rect 2685 189 2731 227
rect 2685 155 2691 189
rect 2725 155 2731 189
rect 2685 117 2731 155
rect 2685 83 2691 117
rect 2725 83 2731 117
rect 2685 45 2731 83
rect 2685 11 2691 45
rect 2725 11 2731 45
rect 2685 -27 2731 11
rect 2685 -61 2691 -27
rect 2725 -61 2731 -27
rect -1881 -181 -1847 -97
rect 235 -143 269 -97
rect 234 -181 269 -143
rect 2351 -181 2385 -97
rect 2685 -100 2731 -61
rect 3743 261 3789 300
rect 3743 227 3749 261
rect 3783 227 3789 261
rect 3743 189 3789 227
rect 3743 155 3749 189
rect 3783 155 3789 189
rect 3743 117 3789 155
rect 3743 83 3749 117
rect 3783 83 3789 117
rect 3743 45 3789 83
rect 3743 11 3749 45
rect 3783 11 3789 45
rect 3743 -27 3789 11
rect 3743 -61 3749 -27
rect 3783 -61 3789 -27
rect 3743 -100 3789 -61
rect 4801 261 4847 300
rect 4801 227 4807 261
rect 4841 227 4847 261
rect 4801 189 4847 227
rect 4801 155 4807 189
rect 4841 155 4847 189
rect 4801 117 4847 155
rect 4801 83 4807 117
rect 4841 83 4847 117
rect 4801 45 4847 83
rect 4801 11 4807 45
rect 4841 11 4847 45
rect 4801 -27 4847 11
rect 4801 -61 4807 -27
rect 4841 -61 4847 -27
rect 4801 -100 4847 -61
rect 5859 261 5905 300
rect 5859 227 5865 261
rect 5899 227 5905 261
rect 5859 189 5905 227
rect 5859 155 5865 189
rect 5899 155 5905 189
rect 5859 117 5905 155
rect 5859 83 5865 117
rect 5899 83 5905 117
rect 5859 45 5905 83
rect 5859 11 5865 45
rect 5899 11 5905 45
rect 5859 -27 5905 11
rect 5859 -61 5865 -27
rect 5899 -61 5905 -27
rect 5859 -100 5905 -61
rect 6917 261 6963 300
rect 6917 227 6923 261
rect 6957 227 6963 261
rect 6917 189 6963 227
rect 6917 155 6923 189
rect 6957 155 6963 189
rect 6917 117 6963 155
rect 6917 83 6923 117
rect 6957 83 6963 117
rect 6917 45 6963 83
rect 6917 11 6923 45
rect 6957 11 6963 45
rect 6917 -27 6963 11
rect 6917 -61 6923 -27
rect 6957 -61 6963 -27
rect 6917 -100 6963 -61
rect 7975 261 8021 300
rect 7975 227 7981 261
rect 8015 227 8021 261
rect 7975 189 8021 227
rect 7975 155 7981 189
rect 8015 155 8021 189
rect 7975 117 8021 155
rect 7975 83 7981 117
rect 8015 83 8021 117
rect 7975 45 8021 83
rect 7975 11 7981 45
rect 8015 11 8021 45
rect 7975 -27 8021 11
rect 7975 -61 7981 -27
rect 8015 -61 8021 -27
rect 7975 -100 8021 -61
rect 3749 -166 3783 -100
rect 5865 -128 5899 -100
rect 5864 -166 5899 -128
rect 7981 -166 8015 -100
rect -1882 -184 2385 -181
rect 3748 -169 8015 -166
rect -1882 -218 2384 -184
rect 3748 -203 8014 -169
rect 2254 -297 2384 -218
rect 3750 -297 4005 -203
rect 2252 -298 4006 -297
rect 2252 -445 4007 -298
use sky130_fd_pr__pfet_g5v0d10v5_9HRSSM  sky130_fd_pr__pfet_g5v0d10v5_9HRSSM_4
timestamp 1640969486
transform 1 0 -2393 0 1 85
box -624 -266 624 266
use sky130_fd_pr__pfet_g5v0d10v5_9HRSSM  sky130_fd_pr__pfet_g5v0d10v5_9HRSSM_3
timestamp 1640969486
transform 1 0 -1335 0 1 85
box -624 -266 624 266
use sky130_fd_pr__pfet_g5v0d10v5_9HRSSM  sky130_fd_pr__pfet_g5v0d10v5_9HRSSM_2
timestamp 1640969486
transform 1 0 -277 0 1 85
box -624 -266 624 266
use sky130_fd_pr__pfet_g5v0d10v5_9HRSSM  sky130_fd_pr__pfet_g5v0d10v5_9HRSSM_1
timestamp 1640969486
transform 1 0 781 0 1 85
box -624 -266 624 266
use sky130_fd_pr__pfet_g5v0d10v5_9HRSSM  sky130_fd_pr__pfet_g5v0d10v5_9HRSSM_0
timestamp 1640969486
transform 1 0 1839 0 1 85
box -624 -266 624 266
<< labels >>
flabel locali s -2619 -207 -2619 -207 0 FreeSans 2500 0 0 0 S
port 1 nsew
flabel locali s 3011 -192 3011 -192 0 FreeSans 2500 0 0 0 S
port 1 nsew
flabel metal1 s 1786 -207 1786 -207 0 FreeSans 2500 0 0 0 D
port 2 nsew
flabel metal1 s 7416 -192 7416 -192 0 FreeSans 2500 0 0 0 D
port 2 nsew
flabel locali s 35 434 35 434 0 FreeSans 2500 0 0 0 G
port 3 nsew
flabel locali s 5665 449 5665 449 0 FreeSans 2500 0 0 0 G
port 3 nsew
<< end >>
