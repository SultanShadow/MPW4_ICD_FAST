magic
tech sky130A
magscale 1 2
timestamp 1640969486
<< pwell >>
rect -191 1302 191 1388
rect -191 -1302 -105 1302
rect 105 -1302 191 1302
rect -191 -1388 191 -1302
<< psubdiff >>
rect -165 1328 -51 1362
rect -17 1328 17 1362
rect 51 1328 165 1362
rect -165 1241 -131 1328
rect 131 1241 165 1328
rect -165 1173 -131 1207
rect -165 1105 -131 1139
rect -165 1037 -131 1071
rect -165 969 -131 1003
rect -165 901 -131 935
rect -165 833 -131 867
rect -165 765 -131 799
rect -165 697 -131 731
rect -165 629 -131 663
rect -165 561 -131 595
rect -165 493 -131 527
rect -165 425 -131 459
rect -165 357 -131 391
rect -165 289 -131 323
rect -165 221 -131 255
rect -165 153 -131 187
rect -165 85 -131 119
rect -165 17 -131 51
rect -165 -51 -131 -17
rect -165 -119 -131 -85
rect -165 -187 -131 -153
rect -165 -255 -131 -221
rect -165 -323 -131 -289
rect -165 -391 -131 -357
rect -165 -459 -131 -425
rect -165 -527 -131 -493
rect -165 -595 -131 -561
rect -165 -663 -131 -629
rect -165 -731 -131 -697
rect -165 -799 -131 -765
rect -165 -867 -131 -833
rect -165 -935 -131 -901
rect -165 -1003 -131 -969
rect -165 -1071 -131 -1037
rect -165 -1139 -131 -1105
rect -165 -1207 -131 -1173
rect 131 1173 165 1207
rect 131 1105 165 1139
rect 131 1037 165 1071
rect 131 969 165 1003
rect 131 901 165 935
rect 131 833 165 867
rect 131 765 165 799
rect 131 697 165 731
rect 131 629 165 663
rect 131 561 165 595
rect 131 493 165 527
rect 131 425 165 459
rect 131 357 165 391
rect 131 289 165 323
rect 131 221 165 255
rect 131 153 165 187
rect 131 85 165 119
rect 131 17 165 51
rect 131 -51 165 -17
rect 131 -119 165 -85
rect 131 -187 165 -153
rect 131 -255 165 -221
rect 131 -323 165 -289
rect 131 -391 165 -357
rect 131 -459 165 -425
rect 131 -527 165 -493
rect 131 -595 165 -561
rect 131 -663 165 -629
rect 131 -731 165 -697
rect 131 -799 165 -765
rect 131 -867 165 -833
rect 131 -935 165 -901
rect 131 -1003 165 -969
rect 131 -1071 165 -1037
rect 131 -1139 165 -1105
rect 131 -1207 165 -1173
rect -165 -1328 -131 -1241
rect 131 -1328 165 -1241
rect -165 -1362 -51 -1328
rect -17 -1362 17 -1328
rect 51 -1362 165 -1328
<< psubdiffcont >>
rect -51 1328 -17 1362
rect 17 1328 51 1362
rect -165 1207 -131 1241
rect -165 1139 -131 1173
rect -165 1071 -131 1105
rect -165 1003 -131 1037
rect -165 935 -131 969
rect -165 867 -131 901
rect -165 799 -131 833
rect -165 731 -131 765
rect -165 663 -131 697
rect -165 595 -131 629
rect -165 527 -131 561
rect -165 459 -131 493
rect -165 391 -131 425
rect -165 323 -131 357
rect -165 255 -131 289
rect -165 187 -131 221
rect -165 119 -131 153
rect -165 51 -131 85
rect -165 -17 -131 17
rect -165 -85 -131 -51
rect -165 -153 -131 -119
rect -165 -221 -131 -187
rect -165 -289 -131 -255
rect -165 -357 -131 -323
rect -165 -425 -131 -391
rect -165 -493 -131 -459
rect -165 -561 -131 -527
rect -165 -629 -131 -595
rect -165 -697 -131 -663
rect -165 -765 -131 -731
rect -165 -833 -131 -799
rect -165 -901 -131 -867
rect -165 -969 -131 -935
rect -165 -1037 -131 -1003
rect -165 -1105 -131 -1071
rect -165 -1173 -131 -1139
rect -165 -1241 -131 -1207
rect 131 1207 165 1241
rect 131 1139 165 1173
rect 131 1071 165 1105
rect 131 1003 165 1037
rect 131 935 165 969
rect 131 867 165 901
rect 131 799 165 833
rect 131 731 165 765
rect 131 663 165 697
rect 131 595 165 629
rect 131 527 165 561
rect 131 459 165 493
rect 131 391 165 425
rect 131 323 165 357
rect 131 255 165 289
rect 131 187 165 221
rect 131 119 165 153
rect 131 51 165 85
rect 131 -17 165 17
rect 131 -85 165 -51
rect 131 -153 165 -119
rect 131 -221 165 -187
rect 131 -289 165 -255
rect 131 -357 165 -323
rect 131 -425 165 -391
rect 131 -493 165 -459
rect 131 -561 165 -527
rect 131 -629 165 -595
rect 131 -697 165 -663
rect 131 -765 165 -731
rect 131 -833 165 -799
rect 131 -901 165 -867
rect 131 -969 165 -935
rect 131 -1037 165 -1003
rect 131 -1105 165 -1071
rect 131 -1173 165 -1139
rect 131 -1241 165 -1207
rect -51 -1362 -17 -1328
rect 17 -1362 51 -1328
<< xpolycontact >>
rect -35 800 35 1232
rect -35 -1232 35 -800
<< ppolyres >>
rect -35 -800 35 800
<< locali >>
rect -165 1328 -51 1362
rect -17 1328 17 1362
rect 51 1328 165 1362
rect -165 1241 -131 1328
rect 131 1241 165 1328
rect -165 1173 -131 1207
rect -165 1105 -131 1139
rect -165 1037 -131 1071
rect -165 969 -131 1003
rect -165 901 -131 935
rect -165 833 -131 867
rect 131 1173 165 1207
rect 131 1105 165 1139
rect 131 1037 165 1071
rect 131 969 165 1003
rect 131 901 165 935
rect 131 833 165 867
rect -165 765 -131 799
rect -165 697 -131 731
rect -165 629 -131 663
rect -165 561 -131 595
rect -165 493 -131 527
rect -165 425 -131 459
rect -165 357 -131 391
rect -165 289 -131 323
rect -165 221 -131 255
rect -165 153 -131 187
rect -165 85 -131 119
rect -165 17 -131 51
rect -165 -51 -131 -17
rect -165 -119 -131 -85
rect -165 -187 -131 -153
rect -165 -255 -131 -221
rect -165 -323 -131 -289
rect -165 -391 -131 -357
rect -165 -459 -131 -425
rect -165 -527 -131 -493
rect -165 -595 -131 -561
rect -165 -663 -131 -629
rect -165 -731 -131 -697
rect -165 -799 -131 -765
rect 131 765 165 799
rect 131 697 165 731
rect 131 629 165 663
rect 131 561 165 595
rect 131 493 165 527
rect 131 425 165 459
rect 131 357 165 391
rect 131 289 165 323
rect 131 221 165 255
rect 131 153 165 187
rect 131 85 165 119
rect 131 17 165 51
rect 131 -51 165 -17
rect 131 -119 165 -85
rect 131 -187 165 -153
rect 131 -255 165 -221
rect 131 -323 165 -289
rect 131 -391 165 -357
rect 131 -459 165 -425
rect 131 -527 165 -493
rect 131 -595 165 -561
rect 131 -663 165 -629
rect 131 -731 165 -697
rect 131 -799 165 -765
rect -165 -867 -131 -833
rect -165 -935 -131 -901
rect -165 -1003 -131 -969
rect -165 -1071 -131 -1037
rect -165 -1139 -131 -1105
rect -165 -1207 -131 -1173
rect 131 -867 165 -833
rect 131 -935 165 -901
rect 131 -1003 165 -969
rect 131 -1071 165 -1037
rect 131 -1139 165 -1105
rect 131 -1207 165 -1173
rect -165 -1328 -131 -1241
rect 131 -1328 165 -1241
rect -165 -1362 -51 -1328
rect -17 -1362 17 -1328
rect 51 -1362 165 -1328
<< viali >>
rect -17 1178 17 1212
rect -17 1106 17 1140
rect -17 1034 17 1068
rect -17 962 17 996
rect -17 890 17 924
rect -17 818 17 852
rect -17 -853 17 -819
rect -17 -925 17 -891
rect -17 -997 17 -963
rect -17 -1069 17 -1035
rect -17 -1141 17 -1107
rect -17 -1213 17 -1179
<< metal1 >>
rect -25 1212 25 1226
rect -25 1178 -17 1212
rect 17 1178 25 1212
rect -25 1140 25 1178
rect -25 1106 -17 1140
rect 17 1106 25 1140
rect -25 1068 25 1106
rect -25 1034 -17 1068
rect 17 1034 25 1068
rect -25 996 25 1034
rect -25 962 -17 996
rect 17 962 25 996
rect -25 924 25 962
rect -25 890 -17 924
rect 17 890 25 924
rect -25 852 25 890
rect -25 818 -17 852
rect 17 818 25 852
rect -25 805 25 818
rect -25 -819 25 -805
rect -25 -853 -17 -819
rect 17 -853 25 -819
rect -25 -891 25 -853
rect -25 -925 -17 -891
rect 17 -925 25 -891
rect -25 -963 25 -925
rect -25 -997 -17 -963
rect 17 -997 25 -963
rect -25 -1035 25 -997
rect -25 -1069 -17 -1035
rect 17 -1069 25 -1035
rect -25 -1107 25 -1069
rect -25 -1141 -17 -1107
rect 17 -1141 25 -1107
rect -25 -1179 25 -1141
rect -25 -1213 -17 -1179
rect 17 -1213 25 -1179
rect -25 -1226 25 -1213
<< properties >>
string FIXED_BBOX -148 -1345 148 1345
<< end >>
