magic
tech sky130A
magscale 1 2
timestamp 1640969486
<< pwell >>
rect -191 637 191 723
rect -191 -637 -105 637
rect 105 -637 191 637
rect -191 -723 191 -637
<< psubdiff >>
rect -165 663 -51 697
rect -17 663 17 697
rect 51 663 165 697
rect -165 595 -131 663
rect 131 595 165 663
rect -165 527 -131 561
rect -165 459 -131 493
rect -165 391 -131 425
rect -165 323 -131 357
rect -165 255 -131 289
rect -165 187 -131 221
rect -165 119 -131 153
rect -165 51 -131 85
rect -165 -17 -131 17
rect -165 -85 -131 -51
rect -165 -153 -131 -119
rect -165 -221 -131 -187
rect -165 -289 -131 -255
rect -165 -357 -131 -323
rect -165 -425 -131 -391
rect -165 -493 -131 -459
rect -165 -561 -131 -527
rect 131 527 165 561
rect 131 459 165 493
rect 131 391 165 425
rect 131 323 165 357
rect 131 255 165 289
rect 131 187 165 221
rect 131 119 165 153
rect 131 51 165 85
rect 131 -17 165 17
rect 131 -85 165 -51
rect 131 -153 165 -119
rect 131 -221 165 -187
rect 131 -289 165 -255
rect 131 -357 165 -323
rect 131 -425 165 -391
rect 131 -493 165 -459
rect 131 -561 165 -527
rect -165 -663 -131 -595
rect 131 -663 165 -595
rect -165 -697 -51 -663
rect -17 -697 17 -663
rect 51 -697 165 -663
<< psubdiffcont >>
rect -51 663 -17 697
rect 17 663 51 697
rect -165 561 -131 595
rect -165 493 -131 527
rect -165 425 -131 459
rect -165 357 -131 391
rect -165 289 -131 323
rect -165 221 -131 255
rect -165 153 -131 187
rect -165 85 -131 119
rect -165 17 -131 51
rect -165 -51 -131 -17
rect -165 -119 -131 -85
rect -165 -187 -131 -153
rect -165 -255 -131 -221
rect -165 -323 -131 -289
rect -165 -391 -131 -357
rect -165 -459 -131 -425
rect -165 -527 -131 -493
rect -165 -595 -131 -561
rect 131 561 165 595
rect 131 493 165 527
rect 131 425 165 459
rect 131 357 165 391
rect 131 289 165 323
rect 131 221 165 255
rect 131 153 165 187
rect 131 85 165 119
rect 131 17 165 51
rect 131 -51 165 -17
rect 131 -119 165 -85
rect 131 -187 165 -153
rect 131 -255 165 -221
rect 131 -323 165 -289
rect 131 -391 165 -357
rect 131 -459 165 -425
rect 131 -527 165 -493
rect 131 -595 165 -561
rect -51 -697 -17 -663
rect 17 -697 51 -663
<< xpolycontact >>
rect -35 135 35 567
rect -35 -567 35 -135
<< xpolyres >>
rect -35 -135 35 135
<< locali >>
rect -165 663 -51 697
rect -17 663 17 697
rect 51 663 165 697
rect -165 595 -131 663
rect 131 595 165 663
rect -165 527 -131 561
rect -165 459 -131 493
rect -165 391 -131 425
rect -165 323 -131 357
rect -165 255 -131 289
rect -165 187 -131 221
rect -165 119 -131 153
rect 131 527 165 561
rect 131 459 165 493
rect 131 391 165 425
rect 131 323 165 357
rect 131 255 165 289
rect 131 187 165 221
rect -165 51 -131 85
rect -165 -17 -131 17
rect -165 -85 -131 -51
rect -165 -153 -131 -119
rect 131 119 165 153
rect 131 51 165 85
rect 131 -17 165 17
rect 131 -85 165 -51
rect -165 -221 -131 -187
rect -165 -289 -131 -255
rect -165 -357 -131 -323
rect -165 -425 -131 -391
rect -165 -493 -131 -459
rect -165 -561 -131 -527
rect 131 -153 165 -119
rect 131 -221 165 -187
rect 131 -289 165 -255
rect 131 -357 165 -323
rect 131 -425 165 -391
rect 131 -493 165 -459
rect 131 -561 165 -527
rect -165 -663 -131 -595
rect 131 -663 165 -595
rect -165 -697 -51 -663
rect -17 -697 17 -663
rect 51 -697 165 -663
<< viali >>
rect -17 513 17 547
rect -17 441 17 475
rect -17 369 17 403
rect -17 297 17 331
rect -17 225 17 259
rect -17 153 17 187
rect -17 -188 17 -154
rect -17 -260 17 -226
rect -17 -332 17 -298
rect -17 -404 17 -370
rect -17 -476 17 -442
rect -17 -548 17 -514
<< metal1 >>
rect -25 547 25 561
rect -25 513 -17 547
rect 17 513 25 547
rect -25 475 25 513
rect -25 441 -17 475
rect 17 441 25 475
rect -25 403 25 441
rect -25 369 -17 403
rect 17 369 25 403
rect -25 331 25 369
rect -25 297 -17 331
rect 17 297 25 331
rect -25 259 25 297
rect -25 225 -17 259
rect 17 225 25 259
rect -25 187 25 225
rect -25 153 -17 187
rect 17 153 25 187
rect -25 140 25 153
rect -25 -154 25 -140
rect -25 -188 -17 -154
rect 17 -188 25 -154
rect -25 -226 25 -188
rect -25 -260 -17 -226
rect 17 -260 25 -226
rect -25 -298 25 -260
rect -25 -332 -17 -298
rect 17 -332 25 -298
rect -25 -370 25 -332
rect -25 -404 -17 -370
rect 17 -404 25 -370
rect -25 -442 25 -404
rect -25 -476 -17 -442
rect 17 -476 25 -442
rect -25 -514 25 -476
rect -25 -548 -17 -514
rect 17 -548 25 -514
rect -25 -561 25 -548
<< properties >>
string FIXED_BBOX -148 -680 148 680
<< end >>
