magic
tech sky130A
magscale 1 2
timestamp 1640969486
<< nwell >>
rect 509 -1491 6581 3083
<< nsubdiff >>
rect 690 2966 6312 2981
rect 690 2660 1709 2966
rect 5755 2660 6312 2966
rect 690 2645 6312 2660
rect 690 2359 974 2645
rect 690 -463 713 2359
rect 951 -463 974 2359
rect 690 -847 974 -463
rect 6028 2315 6312 2645
rect 6028 -507 6051 2315
rect 6289 -507 6312 2315
rect 6028 -847 6312 -507
rect 690 -862 6312 -847
rect 690 -1168 1441 -862
rect 5487 -1168 6312 -862
rect 690 -1183 6312 -1168
<< nsubdiffcont >>
rect 1709 2660 5755 2966
rect 713 -463 951 2359
rect 6051 -507 6289 2315
rect 1441 -1168 5487 -862
<< poly >>
rect 1560 2408 5452 2422
rect 1560 2374 1577 2408
rect 1611 2374 1645 2408
rect 1679 2374 1713 2408
rect 1747 2374 1781 2408
rect 1815 2374 1849 2408
rect 1883 2374 1917 2408
rect 1951 2374 1985 2408
rect 2019 2374 2053 2408
rect 2087 2374 2121 2408
rect 2155 2374 2189 2408
rect 2223 2374 2257 2408
rect 2291 2374 2325 2408
rect 2359 2374 2393 2408
rect 2427 2374 2461 2408
rect 2495 2374 2529 2408
rect 2563 2374 2597 2408
rect 2631 2374 2665 2408
rect 2699 2374 2733 2408
rect 2767 2374 2801 2408
rect 2835 2374 2869 2408
rect 2903 2374 2937 2408
rect 2971 2374 3005 2408
rect 3039 2374 3073 2408
rect 3107 2374 3141 2408
rect 3175 2374 3209 2408
rect 3243 2374 3277 2408
rect 3311 2374 3345 2408
rect 3379 2374 3413 2408
rect 3447 2374 3481 2408
rect 3515 2374 3549 2408
rect 3583 2374 3617 2408
rect 3651 2374 3685 2408
rect 3719 2374 3753 2408
rect 3787 2374 3821 2408
rect 3855 2374 3889 2408
rect 3923 2374 3957 2408
rect 3991 2374 4025 2408
rect 4059 2374 4093 2408
rect 4127 2374 4161 2408
rect 4195 2374 4229 2408
rect 4263 2374 4297 2408
rect 4331 2374 4365 2408
rect 4399 2374 4433 2408
rect 4467 2374 4501 2408
rect 4535 2374 4569 2408
rect 4603 2374 4637 2408
rect 4671 2374 4705 2408
rect 4739 2374 4773 2408
rect 4807 2374 4841 2408
rect 4875 2374 4909 2408
rect 4943 2374 4977 2408
rect 5011 2374 5045 2408
rect 5079 2374 5113 2408
rect 5147 2374 5181 2408
rect 5215 2374 5249 2408
rect 5283 2374 5317 2408
rect 5351 2374 5385 2408
rect 5419 2374 5452 2408
rect 1560 2358 5452 2374
rect 1560 2316 1660 2358
rect 1718 2316 1818 2358
rect 1876 2316 1976 2358
rect 2034 2316 2134 2358
rect 2192 2316 2292 2358
rect 2350 2316 2450 2358
rect 2508 2316 2608 2358
rect 2666 2316 2766 2358
rect 2824 2316 2924 2358
rect 2982 2316 3082 2358
rect 3140 2316 3240 2358
rect 3298 2316 3398 2358
rect 3456 2316 3556 2358
rect 3614 2316 3714 2358
rect 3772 2316 3872 2358
rect 3930 2316 4030 2358
rect 4088 2316 4188 2358
rect 4246 2316 4346 2358
rect 4404 2316 4504 2358
rect 4562 2316 4662 2358
rect 4720 2316 4820 2358
rect 4878 2316 4978 2358
rect 5036 2316 5136 2358
rect 5194 2316 5294 2358
rect 5352 2316 5452 2358
rect 1560 -618 1660 -576
rect 1718 -618 1818 -576
rect 1876 -618 1976 -576
rect 2034 -618 2134 -576
rect 2192 -618 2292 -576
rect 2350 -618 2450 -576
rect 2508 -618 2608 -576
rect 2666 -618 2766 -576
rect 2824 -618 2924 -576
rect 2982 -618 3082 -576
rect 3140 -618 3240 -576
rect 3298 -618 3398 -576
rect 3456 -618 3556 -576
rect 3614 -618 3714 -576
rect 3772 -618 3872 -576
rect 3930 -618 4030 -576
rect 4088 -618 4188 -576
rect 4246 -618 4346 -576
rect 4404 -618 4504 -576
rect 4562 -618 4662 -576
rect 4720 -618 4820 -576
rect 4878 -618 4978 -576
rect 5036 -618 5136 -576
rect 5194 -618 5294 -576
rect 5352 -618 5452 -576
rect 1560 -632 5452 -618
rect 1560 -666 1577 -632
rect 1611 -666 1645 -632
rect 1679 -666 1713 -632
rect 1747 -666 1781 -632
rect 1815 -666 1849 -632
rect 1883 -666 1917 -632
rect 1951 -666 1985 -632
rect 2019 -666 2053 -632
rect 2087 -666 2121 -632
rect 2155 -666 2189 -632
rect 2223 -666 2257 -632
rect 2291 -666 2325 -632
rect 2359 -666 2393 -632
rect 2427 -666 2461 -632
rect 2495 -666 2529 -632
rect 2563 -666 2597 -632
rect 2631 -666 2665 -632
rect 2699 -666 2733 -632
rect 2767 -666 2801 -632
rect 2835 -666 2869 -632
rect 2903 -666 2937 -632
rect 2971 -666 3005 -632
rect 3039 -666 3073 -632
rect 3107 -666 3141 -632
rect 3175 -666 3209 -632
rect 3243 -666 3277 -632
rect 3311 -666 3345 -632
rect 3379 -666 3413 -632
rect 3447 -666 3481 -632
rect 3515 -666 3549 -632
rect 3583 -666 3617 -632
rect 3651 -666 3685 -632
rect 3719 -666 3753 -632
rect 3787 -666 3821 -632
rect 3855 -666 3889 -632
rect 3923 -666 3957 -632
rect 3991 -666 4025 -632
rect 4059 -666 4093 -632
rect 4127 -666 4161 -632
rect 4195 -666 4229 -632
rect 4263 -666 4297 -632
rect 4331 -666 4365 -632
rect 4399 -666 4433 -632
rect 4467 -666 4501 -632
rect 4535 -666 4569 -632
rect 4603 -666 4637 -632
rect 4671 -666 4705 -632
rect 4739 -666 4773 -632
rect 4807 -666 4841 -632
rect 4875 -666 4909 -632
rect 4943 -666 4977 -632
rect 5011 -666 5045 -632
rect 5079 -666 5113 -632
rect 5147 -666 5181 -632
rect 5215 -666 5249 -632
rect 5283 -666 5317 -632
rect 5351 -666 5385 -632
rect 5419 -666 5452 -632
rect 1560 -682 5452 -666
<< polycont >>
rect 1577 2374 1611 2408
rect 1645 2374 1679 2408
rect 1713 2374 1747 2408
rect 1781 2374 1815 2408
rect 1849 2374 1883 2408
rect 1917 2374 1951 2408
rect 1985 2374 2019 2408
rect 2053 2374 2087 2408
rect 2121 2374 2155 2408
rect 2189 2374 2223 2408
rect 2257 2374 2291 2408
rect 2325 2374 2359 2408
rect 2393 2374 2427 2408
rect 2461 2374 2495 2408
rect 2529 2374 2563 2408
rect 2597 2374 2631 2408
rect 2665 2374 2699 2408
rect 2733 2374 2767 2408
rect 2801 2374 2835 2408
rect 2869 2374 2903 2408
rect 2937 2374 2971 2408
rect 3005 2374 3039 2408
rect 3073 2374 3107 2408
rect 3141 2374 3175 2408
rect 3209 2374 3243 2408
rect 3277 2374 3311 2408
rect 3345 2374 3379 2408
rect 3413 2374 3447 2408
rect 3481 2374 3515 2408
rect 3549 2374 3583 2408
rect 3617 2374 3651 2408
rect 3685 2374 3719 2408
rect 3753 2374 3787 2408
rect 3821 2374 3855 2408
rect 3889 2374 3923 2408
rect 3957 2374 3991 2408
rect 4025 2374 4059 2408
rect 4093 2374 4127 2408
rect 4161 2374 4195 2408
rect 4229 2374 4263 2408
rect 4297 2374 4331 2408
rect 4365 2374 4399 2408
rect 4433 2374 4467 2408
rect 4501 2374 4535 2408
rect 4569 2374 4603 2408
rect 4637 2374 4671 2408
rect 4705 2374 4739 2408
rect 4773 2374 4807 2408
rect 4841 2374 4875 2408
rect 4909 2374 4943 2408
rect 4977 2374 5011 2408
rect 5045 2374 5079 2408
rect 5113 2374 5147 2408
rect 5181 2374 5215 2408
rect 5249 2374 5283 2408
rect 5317 2374 5351 2408
rect 5385 2374 5419 2408
rect 1577 -666 1611 -632
rect 1645 -666 1679 -632
rect 1713 -666 1747 -632
rect 1781 -666 1815 -632
rect 1849 -666 1883 -632
rect 1917 -666 1951 -632
rect 1985 -666 2019 -632
rect 2053 -666 2087 -632
rect 2121 -666 2155 -632
rect 2189 -666 2223 -632
rect 2257 -666 2291 -632
rect 2325 -666 2359 -632
rect 2393 -666 2427 -632
rect 2461 -666 2495 -632
rect 2529 -666 2563 -632
rect 2597 -666 2631 -632
rect 2665 -666 2699 -632
rect 2733 -666 2767 -632
rect 2801 -666 2835 -632
rect 2869 -666 2903 -632
rect 2937 -666 2971 -632
rect 3005 -666 3039 -632
rect 3073 -666 3107 -632
rect 3141 -666 3175 -632
rect 3209 -666 3243 -632
rect 3277 -666 3311 -632
rect 3345 -666 3379 -632
rect 3413 -666 3447 -632
rect 3481 -666 3515 -632
rect 3549 -666 3583 -632
rect 3617 -666 3651 -632
rect 3685 -666 3719 -632
rect 3753 -666 3787 -632
rect 3821 -666 3855 -632
rect 3889 -666 3923 -632
rect 3957 -666 3991 -632
rect 4025 -666 4059 -632
rect 4093 -666 4127 -632
rect 4161 -666 4195 -632
rect 4229 -666 4263 -632
rect 4297 -666 4331 -632
rect 4365 -666 4399 -632
rect 4433 -666 4467 -632
rect 4501 -666 4535 -632
rect 4569 -666 4603 -632
rect 4637 -666 4671 -632
rect 4705 -666 4739 -632
rect 4773 -666 4807 -632
rect 4841 -666 4875 -632
rect 4909 -666 4943 -632
rect 4977 -666 5011 -632
rect 5045 -666 5079 -632
rect 5113 -666 5147 -632
rect 5181 -666 5215 -632
rect 5249 -666 5283 -632
rect 5317 -666 5351 -632
rect 5385 -666 5419 -632
<< locali >>
rect 690 2966 6312 2981
rect 690 2660 1709 2966
rect 5755 2660 6312 2966
rect 690 2645 6312 2660
rect 690 2359 974 2645
rect 690 -463 713 2359
rect 951 -463 974 2359
rect 1560 2408 5452 2422
rect 1560 2374 1577 2408
rect 1643 2374 1645 2408
rect 1679 2374 1681 2408
rect 1747 2374 1753 2408
rect 1815 2374 1825 2408
rect 1883 2374 1897 2408
rect 1951 2374 1969 2408
rect 2019 2374 2041 2408
rect 2087 2374 2113 2408
rect 2155 2374 2185 2408
rect 2223 2374 2257 2408
rect 2291 2374 2325 2408
rect 2363 2374 2393 2408
rect 2435 2374 2461 2408
rect 2507 2374 2529 2408
rect 2579 2374 2597 2408
rect 2651 2374 2665 2408
rect 2723 2374 2733 2408
rect 2795 2374 2801 2408
rect 2867 2374 2869 2408
rect 2903 2374 2905 2408
rect 2971 2374 2977 2408
rect 3039 2374 3049 2408
rect 3107 2374 3121 2408
rect 3175 2374 3193 2408
rect 3243 2374 3265 2408
rect 3311 2374 3337 2408
rect 3379 2374 3409 2408
rect 3447 2374 3481 2408
rect 3515 2374 3549 2408
rect 3587 2374 3617 2408
rect 3659 2374 3685 2408
rect 3731 2374 3753 2408
rect 3803 2374 3821 2408
rect 3875 2374 3889 2408
rect 3947 2374 3957 2408
rect 4019 2374 4025 2408
rect 4091 2374 4093 2408
rect 4127 2374 4129 2408
rect 4195 2374 4201 2408
rect 4263 2374 4273 2408
rect 4331 2374 4345 2408
rect 4399 2374 4417 2408
rect 4467 2374 4489 2408
rect 4535 2374 4561 2408
rect 4603 2374 4633 2408
rect 4671 2374 4705 2408
rect 4739 2374 4773 2408
rect 4811 2374 4841 2408
rect 4883 2374 4909 2408
rect 4955 2374 4977 2408
rect 5027 2374 5045 2408
rect 5099 2374 5113 2408
rect 5171 2374 5181 2408
rect 5243 2374 5249 2408
rect 5315 2374 5317 2408
rect 5351 2374 5353 2408
rect 5419 2374 5452 2408
rect 1560 2358 5452 2374
rect 690 -847 974 -463
rect 6028 2315 6312 2645
rect 6028 -507 6051 2315
rect 6289 -507 6312 2315
rect 1560 -632 5452 -618
rect 1560 -666 1577 -632
rect 1643 -666 1645 -632
rect 1679 -666 1681 -632
rect 1747 -666 1753 -632
rect 1815 -666 1825 -632
rect 1883 -666 1897 -632
rect 1951 -666 1969 -632
rect 2019 -666 2041 -632
rect 2087 -666 2113 -632
rect 2155 -666 2185 -632
rect 2223 -666 2257 -632
rect 2291 -666 2325 -632
rect 2363 -666 2393 -632
rect 2435 -666 2461 -632
rect 2507 -666 2529 -632
rect 2579 -666 2597 -632
rect 2651 -666 2665 -632
rect 2723 -666 2733 -632
rect 2795 -666 2801 -632
rect 2867 -666 2869 -632
rect 2903 -666 2905 -632
rect 2971 -666 2977 -632
rect 3039 -666 3049 -632
rect 3107 -666 3121 -632
rect 3175 -666 3193 -632
rect 3243 -666 3265 -632
rect 3311 -666 3337 -632
rect 3379 -666 3409 -632
rect 3447 -666 3481 -632
rect 3515 -666 3549 -632
rect 3587 -666 3617 -632
rect 3659 -666 3685 -632
rect 3731 -666 3753 -632
rect 3803 -666 3821 -632
rect 3875 -666 3889 -632
rect 3947 -666 3957 -632
rect 4019 -666 4025 -632
rect 4091 -666 4093 -632
rect 4127 -666 4129 -632
rect 4195 -666 4201 -632
rect 4263 -666 4273 -632
rect 4331 -666 4345 -632
rect 4399 -666 4417 -632
rect 4467 -666 4489 -632
rect 4535 -666 4561 -632
rect 4603 -666 4633 -632
rect 4671 -666 4705 -632
rect 4739 -666 4773 -632
rect 4811 -666 4841 -632
rect 4883 -666 4909 -632
rect 4955 -666 4977 -632
rect 5027 -666 5045 -632
rect 5099 -666 5113 -632
rect 5171 -666 5181 -632
rect 5243 -666 5249 -632
rect 5315 -666 5317 -632
rect 5351 -666 5353 -632
rect 5419 -666 5452 -632
rect 1560 -682 5452 -666
rect 6028 -847 6312 -507
rect 690 -862 6312 -847
rect 690 -1168 1441 -862
rect 5487 -1168 6312 -862
rect 690 -1183 6312 -1168
<< viali >>
rect 745 1566 923 2176
rect 1609 2374 1611 2408
rect 1611 2374 1643 2408
rect 1681 2374 1713 2408
rect 1713 2374 1715 2408
rect 1753 2374 1781 2408
rect 1781 2374 1787 2408
rect 1825 2374 1849 2408
rect 1849 2374 1859 2408
rect 1897 2374 1917 2408
rect 1917 2374 1931 2408
rect 1969 2374 1985 2408
rect 1985 2374 2003 2408
rect 2041 2374 2053 2408
rect 2053 2374 2075 2408
rect 2113 2374 2121 2408
rect 2121 2374 2147 2408
rect 2185 2374 2189 2408
rect 2189 2374 2219 2408
rect 2257 2374 2291 2408
rect 2329 2374 2359 2408
rect 2359 2374 2363 2408
rect 2401 2374 2427 2408
rect 2427 2374 2435 2408
rect 2473 2374 2495 2408
rect 2495 2374 2507 2408
rect 2545 2374 2563 2408
rect 2563 2374 2579 2408
rect 2617 2374 2631 2408
rect 2631 2374 2651 2408
rect 2689 2374 2699 2408
rect 2699 2374 2723 2408
rect 2761 2374 2767 2408
rect 2767 2374 2795 2408
rect 2833 2374 2835 2408
rect 2835 2374 2867 2408
rect 2905 2374 2937 2408
rect 2937 2374 2939 2408
rect 2977 2374 3005 2408
rect 3005 2374 3011 2408
rect 3049 2374 3073 2408
rect 3073 2374 3083 2408
rect 3121 2374 3141 2408
rect 3141 2374 3155 2408
rect 3193 2374 3209 2408
rect 3209 2374 3227 2408
rect 3265 2374 3277 2408
rect 3277 2374 3299 2408
rect 3337 2374 3345 2408
rect 3345 2374 3371 2408
rect 3409 2374 3413 2408
rect 3413 2374 3443 2408
rect 3481 2374 3515 2408
rect 3553 2374 3583 2408
rect 3583 2374 3587 2408
rect 3625 2374 3651 2408
rect 3651 2374 3659 2408
rect 3697 2374 3719 2408
rect 3719 2374 3731 2408
rect 3769 2374 3787 2408
rect 3787 2374 3803 2408
rect 3841 2374 3855 2408
rect 3855 2374 3875 2408
rect 3913 2374 3923 2408
rect 3923 2374 3947 2408
rect 3985 2374 3991 2408
rect 3991 2374 4019 2408
rect 4057 2374 4059 2408
rect 4059 2374 4091 2408
rect 4129 2374 4161 2408
rect 4161 2374 4163 2408
rect 4201 2374 4229 2408
rect 4229 2374 4235 2408
rect 4273 2374 4297 2408
rect 4297 2374 4307 2408
rect 4345 2374 4365 2408
rect 4365 2374 4379 2408
rect 4417 2374 4433 2408
rect 4433 2374 4451 2408
rect 4489 2374 4501 2408
rect 4501 2374 4523 2408
rect 4561 2374 4569 2408
rect 4569 2374 4595 2408
rect 4633 2374 4637 2408
rect 4637 2374 4667 2408
rect 4705 2374 4739 2408
rect 4777 2374 4807 2408
rect 4807 2374 4811 2408
rect 4849 2374 4875 2408
rect 4875 2374 4883 2408
rect 4921 2374 4943 2408
rect 4943 2374 4955 2408
rect 4993 2374 5011 2408
rect 5011 2374 5027 2408
rect 5065 2374 5079 2408
rect 5079 2374 5099 2408
rect 5137 2374 5147 2408
rect 5147 2374 5171 2408
rect 5209 2374 5215 2408
rect 5215 2374 5243 2408
rect 5281 2374 5283 2408
rect 5283 2374 5315 2408
rect 5353 2374 5385 2408
rect 5385 2374 5387 2408
rect 6082 1577 6260 2187
rect 1609 -666 1611 -632
rect 1611 -666 1643 -632
rect 1681 -666 1713 -632
rect 1713 -666 1715 -632
rect 1753 -666 1781 -632
rect 1781 -666 1787 -632
rect 1825 -666 1849 -632
rect 1849 -666 1859 -632
rect 1897 -666 1917 -632
rect 1917 -666 1931 -632
rect 1969 -666 1985 -632
rect 1985 -666 2003 -632
rect 2041 -666 2053 -632
rect 2053 -666 2075 -632
rect 2113 -666 2121 -632
rect 2121 -666 2147 -632
rect 2185 -666 2189 -632
rect 2189 -666 2219 -632
rect 2257 -666 2291 -632
rect 2329 -666 2359 -632
rect 2359 -666 2363 -632
rect 2401 -666 2427 -632
rect 2427 -666 2435 -632
rect 2473 -666 2495 -632
rect 2495 -666 2507 -632
rect 2545 -666 2563 -632
rect 2563 -666 2579 -632
rect 2617 -666 2631 -632
rect 2631 -666 2651 -632
rect 2689 -666 2699 -632
rect 2699 -666 2723 -632
rect 2761 -666 2767 -632
rect 2767 -666 2795 -632
rect 2833 -666 2835 -632
rect 2835 -666 2867 -632
rect 2905 -666 2937 -632
rect 2937 -666 2939 -632
rect 2977 -666 3005 -632
rect 3005 -666 3011 -632
rect 3049 -666 3073 -632
rect 3073 -666 3083 -632
rect 3121 -666 3141 -632
rect 3141 -666 3155 -632
rect 3193 -666 3209 -632
rect 3209 -666 3227 -632
rect 3265 -666 3277 -632
rect 3277 -666 3299 -632
rect 3337 -666 3345 -632
rect 3345 -666 3371 -632
rect 3409 -666 3413 -632
rect 3413 -666 3443 -632
rect 3481 -666 3515 -632
rect 3553 -666 3583 -632
rect 3583 -666 3587 -632
rect 3625 -666 3651 -632
rect 3651 -666 3659 -632
rect 3697 -666 3719 -632
rect 3719 -666 3731 -632
rect 3769 -666 3787 -632
rect 3787 -666 3803 -632
rect 3841 -666 3855 -632
rect 3855 -666 3875 -632
rect 3913 -666 3923 -632
rect 3923 -666 3947 -632
rect 3985 -666 3991 -632
rect 3991 -666 4019 -632
rect 4057 -666 4059 -632
rect 4059 -666 4091 -632
rect 4129 -666 4161 -632
rect 4161 -666 4163 -632
rect 4201 -666 4229 -632
rect 4229 -666 4235 -632
rect 4273 -666 4297 -632
rect 4297 -666 4307 -632
rect 4345 -666 4365 -632
rect 4365 -666 4379 -632
rect 4417 -666 4433 -632
rect 4433 -666 4451 -632
rect 4489 -666 4501 -632
rect 4501 -666 4523 -632
rect 4561 -666 4569 -632
rect 4569 -666 4595 -632
rect 4633 -666 4637 -632
rect 4637 -666 4667 -632
rect 4705 -666 4739 -632
rect 4777 -666 4807 -632
rect 4807 -666 4811 -632
rect 4849 -666 4875 -632
rect 4875 -666 4883 -632
rect 4921 -666 4943 -632
rect 4943 -666 4955 -632
rect 4993 -666 5011 -632
rect 5011 -666 5027 -632
rect 5065 -666 5079 -632
rect 5079 -666 5099 -632
rect 5137 -666 5147 -632
rect 5147 -666 5171 -632
rect 5209 -666 5215 -632
rect 5215 -666 5243 -632
rect 5281 -666 5283 -632
rect 5283 -666 5315 -632
rect 5353 -666 5385 -632
rect 5385 -666 5387 -632
<< metal1 >>
rect 1265 2408 5731 2422
rect 1265 2374 1609 2408
rect 1643 2374 1681 2408
rect 1715 2374 1753 2408
rect 1787 2374 1825 2408
rect 1859 2374 1897 2408
rect 1931 2374 1969 2408
rect 2003 2374 2041 2408
rect 2075 2374 2113 2408
rect 2147 2374 2185 2408
rect 2219 2374 2257 2408
rect 2291 2374 2329 2408
rect 2363 2374 2401 2408
rect 2435 2374 2473 2408
rect 2507 2374 2545 2408
rect 2579 2374 2617 2408
rect 2651 2374 2689 2408
rect 2723 2374 2761 2408
rect 2795 2374 2833 2408
rect 2867 2374 2905 2408
rect 2939 2374 2977 2408
rect 3011 2374 3049 2408
rect 3083 2374 3121 2408
rect 3155 2374 3193 2408
rect 3227 2374 3265 2408
rect 3299 2374 3337 2408
rect 3371 2374 3409 2408
rect 3443 2374 3481 2408
rect 3515 2374 3553 2408
rect 3587 2374 3625 2408
rect 3659 2374 3697 2408
rect 3731 2374 3769 2408
rect 3803 2374 3841 2408
rect 3875 2374 3913 2408
rect 3947 2374 3985 2408
rect 4019 2374 4057 2408
rect 4091 2374 4129 2408
rect 4163 2374 4201 2408
rect 4235 2374 4273 2408
rect 4307 2374 4345 2408
rect 4379 2374 4417 2408
rect 4451 2374 4489 2408
rect 4523 2374 4561 2408
rect 4595 2374 4633 2408
rect 4667 2374 4705 2408
rect 4739 2374 4777 2408
rect 4811 2374 4849 2408
rect 4883 2374 4921 2408
rect 4955 2374 4993 2408
rect 5027 2374 5065 2408
rect 5099 2374 5137 2408
rect 5171 2374 5209 2408
rect 5243 2374 5281 2408
rect 5315 2374 5353 2408
rect 5387 2374 5731 2408
rect 1265 2358 5731 2374
rect 690 2185 974 2260
rect 690 1557 744 2185
rect 924 1557 974 2185
rect 690 1507 974 1557
rect 1265 -618 1435 2358
rect 1499 2229 1563 2257
rect 1499 2177 1505 2229
rect 1557 2177 1563 2229
rect 1499 2165 1563 2177
rect 1499 2113 1505 2165
rect 1557 2113 1563 2165
rect 1499 2101 1563 2113
rect 1499 2049 1505 2101
rect 1557 2049 1563 2101
rect 1499 2037 1563 2049
rect 1499 1985 1505 2037
rect 1557 1985 1563 2037
rect 1499 1973 1563 1985
rect 1499 1921 1505 1973
rect 1557 1921 1563 1973
rect 1499 1909 1563 1921
rect 1499 1857 1505 1909
rect 1557 1857 1563 1909
rect 1499 1845 1563 1857
rect 1499 1793 1505 1845
rect 1557 1793 1563 1845
rect 1499 1781 1563 1793
rect 1499 1729 1505 1781
rect 1557 1729 1563 1781
rect 1499 1717 1563 1729
rect 1499 1665 1505 1717
rect 1557 1665 1563 1717
rect 1499 1653 1563 1665
rect 1499 1601 1505 1653
rect 1557 1601 1563 1653
rect 1499 1589 1563 1601
rect 1499 1537 1505 1589
rect 1557 1537 1563 1589
rect 1499 1510 1563 1537
rect 1815 2229 1879 2257
rect 1815 2177 1821 2229
rect 1873 2177 1879 2229
rect 1815 2165 1879 2177
rect 1815 2113 1821 2165
rect 1873 2113 1879 2165
rect 1815 2101 1879 2113
rect 1815 2049 1821 2101
rect 1873 2049 1879 2101
rect 1815 2037 1879 2049
rect 1815 1985 1821 2037
rect 1873 1985 1879 2037
rect 1815 1973 1879 1985
rect 1815 1921 1821 1973
rect 1873 1921 1879 1973
rect 1815 1909 1879 1921
rect 1815 1857 1821 1909
rect 1873 1857 1879 1909
rect 1815 1845 1879 1857
rect 1815 1793 1821 1845
rect 1873 1793 1879 1845
rect 1815 1781 1879 1793
rect 1815 1729 1821 1781
rect 1873 1729 1879 1781
rect 1815 1717 1879 1729
rect 1815 1665 1821 1717
rect 1873 1665 1879 1717
rect 1815 1653 1879 1665
rect 1815 1601 1821 1653
rect 1873 1601 1879 1653
rect 1815 1589 1879 1601
rect 1815 1537 1821 1589
rect 1873 1537 1879 1589
rect 1815 1510 1879 1537
rect 2131 2229 2195 2257
rect 2131 2177 2137 2229
rect 2189 2177 2195 2229
rect 2131 2165 2195 2177
rect 2131 2113 2137 2165
rect 2189 2113 2195 2165
rect 2131 2101 2195 2113
rect 2131 2049 2137 2101
rect 2189 2049 2195 2101
rect 2131 2037 2195 2049
rect 2131 1985 2137 2037
rect 2189 1985 2195 2037
rect 2131 1973 2195 1985
rect 2131 1921 2137 1973
rect 2189 1921 2195 1973
rect 2131 1909 2195 1921
rect 2131 1857 2137 1909
rect 2189 1857 2195 1909
rect 2131 1845 2195 1857
rect 2131 1793 2137 1845
rect 2189 1793 2195 1845
rect 2131 1781 2195 1793
rect 2131 1729 2137 1781
rect 2189 1729 2195 1781
rect 2131 1717 2195 1729
rect 2131 1665 2137 1717
rect 2189 1665 2195 1717
rect 2131 1653 2195 1665
rect 2131 1601 2137 1653
rect 2189 1601 2195 1653
rect 2131 1589 2195 1601
rect 2131 1537 2137 1589
rect 2189 1537 2195 1589
rect 2131 1510 2195 1537
rect 2447 2229 2511 2257
rect 2447 2177 2453 2229
rect 2505 2177 2511 2229
rect 2447 2165 2511 2177
rect 2447 2113 2453 2165
rect 2505 2113 2511 2165
rect 2447 2101 2511 2113
rect 2447 2049 2453 2101
rect 2505 2049 2511 2101
rect 2447 2037 2511 2049
rect 2447 1985 2453 2037
rect 2505 1985 2511 2037
rect 2447 1973 2511 1985
rect 2447 1921 2453 1973
rect 2505 1921 2511 1973
rect 2447 1909 2511 1921
rect 2447 1857 2453 1909
rect 2505 1857 2511 1909
rect 2447 1845 2511 1857
rect 2447 1793 2453 1845
rect 2505 1793 2511 1845
rect 2447 1781 2511 1793
rect 2447 1729 2453 1781
rect 2505 1729 2511 1781
rect 2447 1717 2511 1729
rect 2447 1665 2453 1717
rect 2505 1665 2511 1717
rect 2447 1653 2511 1665
rect 2447 1601 2453 1653
rect 2505 1601 2511 1653
rect 2447 1589 2511 1601
rect 2447 1537 2453 1589
rect 2505 1537 2511 1589
rect 2447 1510 2511 1537
rect 2763 2229 2827 2257
rect 2763 2177 2769 2229
rect 2821 2177 2827 2229
rect 2763 2165 2827 2177
rect 2763 2113 2769 2165
rect 2821 2113 2827 2165
rect 2763 2101 2827 2113
rect 2763 2049 2769 2101
rect 2821 2049 2827 2101
rect 2763 2037 2827 2049
rect 2763 1985 2769 2037
rect 2821 1985 2827 2037
rect 2763 1973 2827 1985
rect 2763 1921 2769 1973
rect 2821 1921 2827 1973
rect 2763 1909 2827 1921
rect 2763 1857 2769 1909
rect 2821 1857 2827 1909
rect 2763 1845 2827 1857
rect 2763 1793 2769 1845
rect 2821 1793 2827 1845
rect 2763 1781 2827 1793
rect 2763 1729 2769 1781
rect 2821 1729 2827 1781
rect 2763 1717 2827 1729
rect 2763 1665 2769 1717
rect 2821 1665 2827 1717
rect 2763 1653 2827 1665
rect 2763 1601 2769 1653
rect 2821 1601 2827 1653
rect 2763 1589 2827 1601
rect 2763 1537 2769 1589
rect 2821 1537 2827 1589
rect 2763 1510 2827 1537
rect 3079 2229 3143 2257
rect 3079 2177 3085 2229
rect 3137 2177 3143 2229
rect 3079 2165 3143 2177
rect 3079 2113 3085 2165
rect 3137 2113 3143 2165
rect 3079 2101 3143 2113
rect 3079 2049 3085 2101
rect 3137 2049 3143 2101
rect 3079 2037 3143 2049
rect 3079 1985 3085 2037
rect 3137 1985 3143 2037
rect 3079 1973 3143 1985
rect 3079 1921 3085 1973
rect 3137 1921 3143 1973
rect 3079 1909 3143 1921
rect 3079 1857 3085 1909
rect 3137 1857 3143 1909
rect 3079 1845 3143 1857
rect 3079 1793 3085 1845
rect 3137 1793 3143 1845
rect 3079 1781 3143 1793
rect 3079 1729 3085 1781
rect 3137 1729 3143 1781
rect 3079 1717 3143 1729
rect 3079 1665 3085 1717
rect 3137 1665 3143 1717
rect 3079 1653 3143 1665
rect 3079 1601 3085 1653
rect 3137 1601 3143 1653
rect 3079 1589 3143 1601
rect 3079 1537 3085 1589
rect 3137 1537 3143 1589
rect 3079 1510 3143 1537
rect 3395 2229 3459 2257
rect 3395 2177 3401 2229
rect 3453 2177 3459 2229
rect 3395 2165 3459 2177
rect 3395 2113 3401 2165
rect 3453 2113 3459 2165
rect 3395 2101 3459 2113
rect 3395 2049 3401 2101
rect 3453 2049 3459 2101
rect 3395 2037 3459 2049
rect 3395 1985 3401 2037
rect 3453 1985 3459 2037
rect 3395 1973 3459 1985
rect 3395 1921 3401 1973
rect 3453 1921 3459 1973
rect 3395 1909 3459 1921
rect 3395 1857 3401 1909
rect 3453 1857 3459 1909
rect 3395 1845 3459 1857
rect 3395 1793 3401 1845
rect 3453 1793 3459 1845
rect 3395 1781 3459 1793
rect 3395 1729 3401 1781
rect 3453 1729 3459 1781
rect 3395 1717 3459 1729
rect 3395 1665 3401 1717
rect 3453 1665 3459 1717
rect 3395 1653 3459 1665
rect 3395 1601 3401 1653
rect 3453 1601 3459 1653
rect 3395 1589 3459 1601
rect 3395 1537 3401 1589
rect 3453 1537 3459 1589
rect 3395 1510 3459 1537
rect 3711 2229 3775 2257
rect 3711 2177 3717 2229
rect 3769 2177 3775 2229
rect 3711 2165 3775 2177
rect 3711 2113 3717 2165
rect 3769 2113 3775 2165
rect 3711 2101 3775 2113
rect 3711 2049 3717 2101
rect 3769 2049 3775 2101
rect 3711 2037 3775 2049
rect 3711 1985 3717 2037
rect 3769 1985 3775 2037
rect 3711 1973 3775 1985
rect 3711 1921 3717 1973
rect 3769 1921 3775 1973
rect 3711 1909 3775 1921
rect 3711 1857 3717 1909
rect 3769 1857 3775 1909
rect 3711 1845 3775 1857
rect 3711 1793 3717 1845
rect 3769 1793 3775 1845
rect 3711 1781 3775 1793
rect 3711 1729 3717 1781
rect 3769 1729 3775 1781
rect 3711 1717 3775 1729
rect 3711 1665 3717 1717
rect 3769 1665 3775 1717
rect 3711 1653 3775 1665
rect 3711 1601 3717 1653
rect 3769 1601 3775 1653
rect 3711 1589 3775 1601
rect 3711 1537 3717 1589
rect 3769 1537 3775 1589
rect 3711 1510 3775 1537
rect 4027 2229 4091 2257
rect 4027 2177 4033 2229
rect 4085 2177 4091 2229
rect 4027 2165 4091 2177
rect 4027 2113 4033 2165
rect 4085 2113 4091 2165
rect 4027 2101 4091 2113
rect 4027 2049 4033 2101
rect 4085 2049 4091 2101
rect 4027 2037 4091 2049
rect 4027 1985 4033 2037
rect 4085 1985 4091 2037
rect 4027 1973 4091 1985
rect 4027 1921 4033 1973
rect 4085 1921 4091 1973
rect 4027 1909 4091 1921
rect 4027 1857 4033 1909
rect 4085 1857 4091 1909
rect 4027 1845 4091 1857
rect 4027 1793 4033 1845
rect 4085 1793 4091 1845
rect 4027 1781 4091 1793
rect 4027 1729 4033 1781
rect 4085 1729 4091 1781
rect 4027 1717 4091 1729
rect 4027 1665 4033 1717
rect 4085 1665 4091 1717
rect 4027 1653 4091 1665
rect 4027 1601 4033 1653
rect 4085 1601 4091 1653
rect 4027 1589 4091 1601
rect 4027 1537 4033 1589
rect 4085 1537 4091 1589
rect 4027 1510 4091 1537
rect 4343 2229 4407 2257
rect 4343 2177 4349 2229
rect 4401 2177 4407 2229
rect 4343 2165 4407 2177
rect 4343 2113 4349 2165
rect 4401 2113 4407 2165
rect 4343 2101 4407 2113
rect 4343 2049 4349 2101
rect 4401 2049 4407 2101
rect 4343 2037 4407 2049
rect 4343 1985 4349 2037
rect 4401 1985 4407 2037
rect 4343 1973 4407 1985
rect 4343 1921 4349 1973
rect 4401 1921 4407 1973
rect 4343 1909 4407 1921
rect 4343 1857 4349 1909
rect 4401 1857 4407 1909
rect 4343 1845 4407 1857
rect 4343 1793 4349 1845
rect 4401 1793 4407 1845
rect 4343 1781 4407 1793
rect 4343 1729 4349 1781
rect 4401 1729 4407 1781
rect 4343 1717 4407 1729
rect 4343 1665 4349 1717
rect 4401 1665 4407 1717
rect 4343 1653 4407 1665
rect 4343 1601 4349 1653
rect 4401 1601 4407 1653
rect 4343 1589 4407 1601
rect 4343 1537 4349 1589
rect 4401 1537 4407 1589
rect 4343 1510 4407 1537
rect 4659 2229 4723 2257
rect 4659 2177 4665 2229
rect 4717 2177 4723 2229
rect 4659 2165 4723 2177
rect 4659 2113 4665 2165
rect 4717 2113 4723 2165
rect 4659 2101 4723 2113
rect 4659 2049 4665 2101
rect 4717 2049 4723 2101
rect 4659 2037 4723 2049
rect 4659 1985 4665 2037
rect 4717 1985 4723 2037
rect 4659 1973 4723 1985
rect 4659 1921 4665 1973
rect 4717 1921 4723 1973
rect 4659 1909 4723 1921
rect 4659 1857 4665 1909
rect 4717 1857 4723 1909
rect 4659 1845 4723 1857
rect 4659 1793 4665 1845
rect 4717 1793 4723 1845
rect 4659 1781 4723 1793
rect 4659 1729 4665 1781
rect 4717 1729 4723 1781
rect 4659 1717 4723 1729
rect 4659 1665 4665 1717
rect 4717 1665 4723 1717
rect 4659 1653 4723 1665
rect 4659 1601 4665 1653
rect 4717 1601 4723 1653
rect 4659 1589 4723 1601
rect 4659 1537 4665 1589
rect 4717 1537 4723 1589
rect 4659 1510 4723 1537
rect 4975 2229 5039 2257
rect 4975 2177 4981 2229
rect 5033 2177 5039 2229
rect 4975 2165 5039 2177
rect 4975 2113 4981 2165
rect 5033 2113 5039 2165
rect 4975 2101 5039 2113
rect 4975 2049 4981 2101
rect 5033 2049 5039 2101
rect 4975 2037 5039 2049
rect 4975 1985 4981 2037
rect 5033 1985 5039 2037
rect 4975 1973 5039 1985
rect 4975 1921 4981 1973
rect 5033 1921 5039 1973
rect 4975 1909 5039 1921
rect 4975 1857 4981 1909
rect 5033 1857 5039 1909
rect 4975 1845 5039 1857
rect 4975 1793 4981 1845
rect 5033 1793 5039 1845
rect 4975 1781 5039 1793
rect 4975 1729 4981 1781
rect 5033 1729 5039 1781
rect 4975 1717 5039 1729
rect 4975 1665 4981 1717
rect 5033 1665 5039 1717
rect 4975 1653 5039 1665
rect 4975 1601 4981 1653
rect 5033 1601 5039 1653
rect 4975 1589 5039 1601
rect 4975 1537 4981 1589
rect 5033 1537 5039 1589
rect 4975 1510 5039 1537
rect 5291 2229 5355 2257
rect 5291 2177 5297 2229
rect 5349 2177 5355 2229
rect 5291 2165 5355 2177
rect 5291 2113 5297 2165
rect 5349 2113 5355 2165
rect 5291 2101 5355 2113
rect 5291 2049 5297 2101
rect 5349 2049 5355 2101
rect 5291 2037 5355 2049
rect 5291 1985 5297 2037
rect 5349 1985 5355 2037
rect 5291 1973 5355 1985
rect 5291 1921 5297 1973
rect 5349 1921 5355 1973
rect 5291 1909 5355 1921
rect 5291 1857 5297 1909
rect 5349 1857 5355 1909
rect 5291 1845 5355 1857
rect 5291 1793 5297 1845
rect 5349 1793 5355 1845
rect 5291 1781 5355 1793
rect 5291 1729 5297 1781
rect 5349 1729 5355 1781
rect 5291 1717 5355 1729
rect 5291 1665 5297 1717
rect 5349 1665 5355 1717
rect 5291 1653 5355 1665
rect 5291 1601 5297 1653
rect 5349 1601 5355 1653
rect 5291 1589 5355 1601
rect 5291 1537 5297 1589
rect 5349 1537 5355 1589
rect 5291 1510 5355 1537
rect 1657 390 1721 424
rect 1657 338 1663 390
rect 1715 338 1721 390
rect 1657 326 1721 338
rect 1657 274 1663 326
rect 1715 274 1721 326
rect 1657 262 1721 274
rect 1657 210 1663 262
rect 1715 210 1721 262
rect 1657 198 1721 210
rect 1657 146 1663 198
rect 1715 146 1721 198
rect 1657 134 1721 146
rect 1657 82 1663 134
rect 1715 82 1721 134
rect 1657 70 1721 82
rect 1657 18 1663 70
rect 1715 18 1721 70
rect 1657 6 1721 18
rect 1657 -46 1663 6
rect 1715 -46 1721 6
rect 1657 -58 1721 -46
rect 1657 -110 1663 -58
rect 1715 -110 1721 -58
rect 1657 -122 1721 -110
rect 1657 -174 1663 -122
rect 1715 -174 1721 -122
rect 1657 -186 1721 -174
rect 1657 -238 1663 -186
rect 1715 -238 1721 -186
rect 1657 -250 1721 -238
rect 1657 -302 1663 -250
rect 1715 -302 1721 -250
rect 1657 -327 1721 -302
rect 1973 390 2037 424
rect 1973 338 1979 390
rect 2031 338 2037 390
rect 1973 326 2037 338
rect 1973 274 1979 326
rect 2031 274 2037 326
rect 1973 262 2037 274
rect 1973 210 1979 262
rect 2031 210 2037 262
rect 1973 198 2037 210
rect 1973 146 1979 198
rect 2031 146 2037 198
rect 1973 134 2037 146
rect 1973 82 1979 134
rect 2031 82 2037 134
rect 1973 70 2037 82
rect 1973 18 1979 70
rect 2031 18 2037 70
rect 1973 6 2037 18
rect 1973 -46 1979 6
rect 2031 -46 2037 6
rect 1973 -58 2037 -46
rect 1973 -110 1979 -58
rect 2031 -110 2037 -58
rect 1973 -122 2037 -110
rect 1973 -174 1979 -122
rect 2031 -174 2037 -122
rect 1973 -186 2037 -174
rect 1973 -238 1979 -186
rect 2031 -238 2037 -186
rect 1973 -250 2037 -238
rect 1973 -302 1979 -250
rect 2031 -302 2037 -250
rect 1973 -327 2037 -302
rect 2289 390 2353 424
rect 2289 338 2295 390
rect 2347 338 2353 390
rect 2289 326 2353 338
rect 2289 274 2295 326
rect 2347 274 2353 326
rect 2289 262 2353 274
rect 2289 210 2295 262
rect 2347 210 2353 262
rect 2289 198 2353 210
rect 2289 146 2295 198
rect 2347 146 2353 198
rect 2289 134 2353 146
rect 2289 82 2295 134
rect 2347 82 2353 134
rect 2289 70 2353 82
rect 2289 18 2295 70
rect 2347 18 2353 70
rect 2289 6 2353 18
rect 2289 -46 2295 6
rect 2347 -46 2353 6
rect 2289 -58 2353 -46
rect 2289 -110 2295 -58
rect 2347 -110 2353 -58
rect 2289 -122 2353 -110
rect 2289 -174 2295 -122
rect 2347 -174 2353 -122
rect 2289 -186 2353 -174
rect 2289 -238 2295 -186
rect 2347 -238 2353 -186
rect 2289 -250 2353 -238
rect 2289 -302 2295 -250
rect 2347 -302 2353 -250
rect 2289 -327 2353 -302
rect 2605 390 2669 424
rect 2605 338 2611 390
rect 2663 338 2669 390
rect 2605 326 2669 338
rect 2605 274 2611 326
rect 2663 274 2669 326
rect 2605 262 2669 274
rect 2605 210 2611 262
rect 2663 210 2669 262
rect 2605 198 2669 210
rect 2605 146 2611 198
rect 2663 146 2669 198
rect 2605 134 2669 146
rect 2605 82 2611 134
rect 2663 82 2669 134
rect 2605 70 2669 82
rect 2605 18 2611 70
rect 2663 18 2669 70
rect 2605 6 2669 18
rect 2605 -46 2611 6
rect 2663 -46 2669 6
rect 2605 -58 2669 -46
rect 2605 -110 2611 -58
rect 2663 -110 2669 -58
rect 2605 -122 2669 -110
rect 2605 -174 2611 -122
rect 2663 -174 2669 -122
rect 2605 -186 2669 -174
rect 2605 -238 2611 -186
rect 2663 -238 2669 -186
rect 2605 -250 2669 -238
rect 2605 -302 2611 -250
rect 2663 -302 2669 -250
rect 2605 -327 2669 -302
rect 2921 390 2985 424
rect 2921 338 2927 390
rect 2979 338 2985 390
rect 2921 326 2985 338
rect 2921 274 2927 326
rect 2979 274 2985 326
rect 2921 262 2985 274
rect 2921 210 2927 262
rect 2979 210 2985 262
rect 2921 198 2985 210
rect 2921 146 2927 198
rect 2979 146 2985 198
rect 2921 134 2985 146
rect 2921 82 2927 134
rect 2979 82 2985 134
rect 2921 70 2985 82
rect 2921 18 2927 70
rect 2979 18 2985 70
rect 2921 6 2985 18
rect 2921 -46 2927 6
rect 2979 -46 2985 6
rect 2921 -58 2985 -46
rect 2921 -110 2927 -58
rect 2979 -110 2985 -58
rect 2921 -122 2985 -110
rect 2921 -174 2927 -122
rect 2979 -174 2985 -122
rect 2921 -186 2985 -174
rect 2921 -238 2927 -186
rect 2979 -238 2985 -186
rect 2921 -250 2985 -238
rect 2921 -302 2927 -250
rect 2979 -302 2985 -250
rect 2921 -327 2985 -302
rect 3237 390 3301 424
rect 3237 338 3243 390
rect 3295 338 3301 390
rect 3237 326 3301 338
rect 3237 274 3243 326
rect 3295 274 3301 326
rect 3237 262 3301 274
rect 3237 210 3243 262
rect 3295 210 3301 262
rect 3237 198 3301 210
rect 3237 146 3243 198
rect 3295 146 3301 198
rect 3237 134 3301 146
rect 3237 82 3243 134
rect 3295 82 3301 134
rect 3237 70 3301 82
rect 3237 18 3243 70
rect 3295 18 3301 70
rect 3237 6 3301 18
rect 3237 -46 3243 6
rect 3295 -46 3301 6
rect 3237 -58 3301 -46
rect 3237 -110 3243 -58
rect 3295 -110 3301 -58
rect 3237 -122 3301 -110
rect 3237 -174 3243 -122
rect 3295 -174 3301 -122
rect 3237 -186 3301 -174
rect 3237 -238 3243 -186
rect 3295 -238 3301 -186
rect 3237 -250 3301 -238
rect 3237 -302 3243 -250
rect 3295 -302 3301 -250
rect 3237 -327 3301 -302
rect 3553 390 3617 424
rect 3553 338 3559 390
rect 3611 338 3617 390
rect 3553 326 3617 338
rect 3553 274 3559 326
rect 3611 274 3617 326
rect 3553 262 3617 274
rect 3553 210 3559 262
rect 3611 210 3617 262
rect 3553 198 3617 210
rect 3553 146 3559 198
rect 3611 146 3617 198
rect 3553 134 3617 146
rect 3553 82 3559 134
rect 3611 82 3617 134
rect 3553 70 3617 82
rect 3553 18 3559 70
rect 3611 18 3617 70
rect 3553 6 3617 18
rect 3553 -46 3559 6
rect 3611 -46 3617 6
rect 3553 -58 3617 -46
rect 3553 -110 3559 -58
rect 3611 -110 3617 -58
rect 3553 -122 3617 -110
rect 3553 -174 3559 -122
rect 3611 -174 3617 -122
rect 3553 -186 3617 -174
rect 3553 -238 3559 -186
rect 3611 -238 3617 -186
rect 3553 -250 3617 -238
rect 3553 -302 3559 -250
rect 3611 -302 3617 -250
rect 3553 -327 3617 -302
rect 3869 390 3933 424
rect 3869 338 3875 390
rect 3927 338 3933 390
rect 3869 326 3933 338
rect 3869 274 3875 326
rect 3927 274 3933 326
rect 3869 262 3933 274
rect 3869 210 3875 262
rect 3927 210 3933 262
rect 3869 198 3933 210
rect 3869 146 3875 198
rect 3927 146 3933 198
rect 3869 134 3933 146
rect 3869 82 3875 134
rect 3927 82 3933 134
rect 3869 70 3933 82
rect 3869 18 3875 70
rect 3927 18 3933 70
rect 3869 6 3933 18
rect 3869 -46 3875 6
rect 3927 -46 3933 6
rect 3869 -58 3933 -46
rect 3869 -110 3875 -58
rect 3927 -110 3933 -58
rect 3869 -122 3933 -110
rect 3869 -174 3875 -122
rect 3927 -174 3933 -122
rect 3869 -186 3933 -174
rect 3869 -238 3875 -186
rect 3927 -238 3933 -186
rect 3869 -250 3933 -238
rect 3869 -302 3875 -250
rect 3927 -302 3933 -250
rect 3869 -327 3933 -302
rect 4185 390 4249 424
rect 4185 338 4191 390
rect 4243 338 4249 390
rect 4185 326 4249 338
rect 4185 274 4191 326
rect 4243 274 4249 326
rect 4185 262 4249 274
rect 4185 210 4191 262
rect 4243 210 4249 262
rect 4185 198 4249 210
rect 4185 146 4191 198
rect 4243 146 4249 198
rect 4185 134 4249 146
rect 4185 82 4191 134
rect 4243 82 4249 134
rect 4185 70 4249 82
rect 4185 18 4191 70
rect 4243 18 4249 70
rect 4185 6 4249 18
rect 4185 -46 4191 6
rect 4243 -46 4249 6
rect 4185 -58 4249 -46
rect 4185 -110 4191 -58
rect 4243 -110 4249 -58
rect 4185 -122 4249 -110
rect 4185 -174 4191 -122
rect 4243 -174 4249 -122
rect 4185 -186 4249 -174
rect 4185 -238 4191 -186
rect 4243 -238 4249 -186
rect 4185 -250 4249 -238
rect 4185 -302 4191 -250
rect 4243 -302 4249 -250
rect 4185 -327 4249 -302
rect 4501 390 4565 424
rect 4501 338 4507 390
rect 4559 338 4565 390
rect 4501 326 4565 338
rect 4501 274 4507 326
rect 4559 274 4565 326
rect 4501 262 4565 274
rect 4501 210 4507 262
rect 4559 210 4565 262
rect 4501 198 4565 210
rect 4501 146 4507 198
rect 4559 146 4565 198
rect 4501 134 4565 146
rect 4501 82 4507 134
rect 4559 82 4565 134
rect 4501 70 4565 82
rect 4501 18 4507 70
rect 4559 18 4565 70
rect 4501 6 4565 18
rect 4501 -46 4507 6
rect 4559 -46 4565 6
rect 4501 -58 4565 -46
rect 4501 -110 4507 -58
rect 4559 -110 4565 -58
rect 4501 -122 4565 -110
rect 4501 -174 4507 -122
rect 4559 -174 4565 -122
rect 4501 -186 4565 -174
rect 4501 -238 4507 -186
rect 4559 -238 4565 -186
rect 4501 -250 4565 -238
rect 4501 -302 4507 -250
rect 4559 -302 4565 -250
rect 4501 -327 4565 -302
rect 4817 390 4881 424
rect 4817 338 4823 390
rect 4875 338 4881 390
rect 4817 326 4881 338
rect 4817 274 4823 326
rect 4875 274 4881 326
rect 4817 262 4881 274
rect 4817 210 4823 262
rect 4875 210 4881 262
rect 4817 198 4881 210
rect 4817 146 4823 198
rect 4875 146 4881 198
rect 4817 134 4881 146
rect 4817 82 4823 134
rect 4875 82 4881 134
rect 4817 70 4881 82
rect 4817 18 4823 70
rect 4875 18 4881 70
rect 4817 6 4881 18
rect 4817 -46 4823 6
rect 4875 -46 4881 6
rect 4817 -58 4881 -46
rect 4817 -110 4823 -58
rect 4875 -110 4881 -58
rect 4817 -122 4881 -110
rect 4817 -174 4823 -122
rect 4875 -174 4881 -122
rect 4817 -186 4881 -174
rect 4817 -238 4823 -186
rect 4875 -238 4881 -186
rect 4817 -250 4881 -238
rect 4817 -302 4823 -250
rect 4875 -302 4881 -250
rect 4817 -327 4881 -302
rect 5133 390 5197 424
rect 5133 338 5139 390
rect 5191 338 5197 390
rect 5133 326 5197 338
rect 5133 274 5139 326
rect 5191 274 5197 326
rect 5133 262 5197 274
rect 5133 210 5139 262
rect 5191 210 5197 262
rect 5133 198 5197 210
rect 5133 146 5139 198
rect 5191 146 5197 198
rect 5133 134 5197 146
rect 5133 82 5139 134
rect 5191 82 5197 134
rect 5133 70 5197 82
rect 5133 18 5139 70
rect 5191 18 5197 70
rect 5133 6 5197 18
rect 5133 -46 5139 6
rect 5191 -46 5197 6
rect 5133 -58 5197 -46
rect 5133 -110 5139 -58
rect 5191 -110 5197 -58
rect 5133 -122 5197 -110
rect 5133 -174 5139 -122
rect 5191 -174 5197 -122
rect 5133 -186 5197 -174
rect 5133 -238 5139 -186
rect 5191 -238 5197 -186
rect 5133 -250 5197 -238
rect 5133 -302 5139 -250
rect 5191 -302 5197 -250
rect 5133 -327 5197 -302
rect 5449 390 5513 424
rect 5449 338 5455 390
rect 5507 338 5513 390
rect 5449 326 5513 338
rect 5449 274 5455 326
rect 5507 274 5513 326
rect 5449 262 5513 274
rect 5449 210 5455 262
rect 5507 210 5513 262
rect 5449 198 5513 210
rect 5449 146 5455 198
rect 5507 146 5513 198
rect 5449 134 5513 146
rect 5449 82 5455 134
rect 5507 82 5513 134
rect 5449 70 5513 82
rect 5449 18 5455 70
rect 5507 18 5513 70
rect 5449 6 5513 18
rect 5449 -46 5455 6
rect 5507 -46 5513 6
rect 5449 -58 5513 -46
rect 5449 -110 5455 -58
rect 5507 -110 5513 -58
rect 5449 -122 5513 -110
rect 5449 -174 5455 -122
rect 5507 -174 5513 -122
rect 5449 -186 5513 -174
rect 5449 -238 5455 -186
rect 5507 -238 5513 -186
rect 5449 -250 5513 -238
rect 5449 -302 5455 -250
rect 5507 -302 5513 -250
rect 5449 -327 5513 -302
rect 5561 -618 5731 2358
rect 6028 2196 6312 2260
rect 6028 1568 6081 2196
rect 6261 1568 6312 2196
rect 6028 1507 6312 1568
rect 1265 -632 5731 -618
rect 1265 -666 1609 -632
rect 1643 -666 1681 -632
rect 1715 -666 1753 -632
rect 1787 -666 1825 -632
rect 1859 -666 1897 -632
rect 1931 -666 1969 -632
rect 2003 -666 2041 -632
rect 2075 -666 2113 -632
rect 2147 -666 2185 -632
rect 2219 -666 2257 -632
rect 2291 -666 2329 -632
rect 2363 -666 2401 -632
rect 2435 -666 2473 -632
rect 2507 -666 2545 -632
rect 2579 -666 2617 -632
rect 2651 -666 2689 -632
rect 2723 -666 2761 -632
rect 2795 -666 2833 -632
rect 2867 -666 2905 -632
rect 2939 -666 2977 -632
rect 3011 -666 3049 -632
rect 3083 -666 3121 -632
rect 3155 -666 3193 -632
rect 3227 -666 3265 -632
rect 3299 -666 3337 -632
rect 3371 -666 3409 -632
rect 3443 -666 3481 -632
rect 3515 -666 3553 -632
rect 3587 -666 3625 -632
rect 3659 -666 3697 -632
rect 3731 -666 3769 -632
rect 3803 -666 3841 -632
rect 3875 -666 3913 -632
rect 3947 -666 3985 -632
rect 4019 -666 4057 -632
rect 4091 -666 4129 -632
rect 4163 -666 4201 -632
rect 4235 -666 4273 -632
rect 4307 -666 4345 -632
rect 4379 -666 4417 -632
rect 4451 -666 4489 -632
rect 4523 -666 4561 -632
rect 4595 -666 4633 -632
rect 4667 -666 4705 -632
rect 4739 -666 4777 -632
rect 4811 -666 4849 -632
rect 4883 -666 4921 -632
rect 4955 -666 4993 -632
rect 5027 -666 5065 -632
rect 5099 -666 5137 -632
rect 5171 -666 5209 -632
rect 5243 -666 5281 -632
rect 5315 -666 5353 -632
rect 5387 -666 5731 -632
rect 1265 -682 5731 -666
<< via1 >>
rect 744 2176 924 2185
rect 744 1566 745 2176
rect 745 1566 923 2176
rect 923 1566 924 2176
rect 744 1557 924 1566
rect 1505 2177 1557 2229
rect 1505 2113 1557 2165
rect 1505 2049 1557 2101
rect 1505 1985 1557 2037
rect 1505 1921 1557 1973
rect 1505 1857 1557 1909
rect 1505 1793 1557 1845
rect 1505 1729 1557 1781
rect 1505 1665 1557 1717
rect 1505 1601 1557 1653
rect 1505 1537 1557 1589
rect 1821 2177 1873 2229
rect 1821 2113 1873 2165
rect 1821 2049 1873 2101
rect 1821 1985 1873 2037
rect 1821 1921 1873 1973
rect 1821 1857 1873 1909
rect 1821 1793 1873 1845
rect 1821 1729 1873 1781
rect 1821 1665 1873 1717
rect 1821 1601 1873 1653
rect 1821 1537 1873 1589
rect 2137 2177 2189 2229
rect 2137 2113 2189 2165
rect 2137 2049 2189 2101
rect 2137 1985 2189 2037
rect 2137 1921 2189 1973
rect 2137 1857 2189 1909
rect 2137 1793 2189 1845
rect 2137 1729 2189 1781
rect 2137 1665 2189 1717
rect 2137 1601 2189 1653
rect 2137 1537 2189 1589
rect 2453 2177 2505 2229
rect 2453 2113 2505 2165
rect 2453 2049 2505 2101
rect 2453 1985 2505 2037
rect 2453 1921 2505 1973
rect 2453 1857 2505 1909
rect 2453 1793 2505 1845
rect 2453 1729 2505 1781
rect 2453 1665 2505 1717
rect 2453 1601 2505 1653
rect 2453 1537 2505 1589
rect 2769 2177 2821 2229
rect 2769 2113 2821 2165
rect 2769 2049 2821 2101
rect 2769 1985 2821 2037
rect 2769 1921 2821 1973
rect 2769 1857 2821 1909
rect 2769 1793 2821 1845
rect 2769 1729 2821 1781
rect 2769 1665 2821 1717
rect 2769 1601 2821 1653
rect 2769 1537 2821 1589
rect 3085 2177 3137 2229
rect 3085 2113 3137 2165
rect 3085 2049 3137 2101
rect 3085 1985 3137 2037
rect 3085 1921 3137 1973
rect 3085 1857 3137 1909
rect 3085 1793 3137 1845
rect 3085 1729 3137 1781
rect 3085 1665 3137 1717
rect 3085 1601 3137 1653
rect 3085 1537 3137 1589
rect 3401 2177 3453 2229
rect 3401 2113 3453 2165
rect 3401 2049 3453 2101
rect 3401 1985 3453 2037
rect 3401 1921 3453 1973
rect 3401 1857 3453 1909
rect 3401 1793 3453 1845
rect 3401 1729 3453 1781
rect 3401 1665 3453 1717
rect 3401 1601 3453 1653
rect 3401 1537 3453 1589
rect 3717 2177 3769 2229
rect 3717 2113 3769 2165
rect 3717 2049 3769 2101
rect 3717 1985 3769 2037
rect 3717 1921 3769 1973
rect 3717 1857 3769 1909
rect 3717 1793 3769 1845
rect 3717 1729 3769 1781
rect 3717 1665 3769 1717
rect 3717 1601 3769 1653
rect 3717 1537 3769 1589
rect 4033 2177 4085 2229
rect 4033 2113 4085 2165
rect 4033 2049 4085 2101
rect 4033 1985 4085 2037
rect 4033 1921 4085 1973
rect 4033 1857 4085 1909
rect 4033 1793 4085 1845
rect 4033 1729 4085 1781
rect 4033 1665 4085 1717
rect 4033 1601 4085 1653
rect 4033 1537 4085 1589
rect 4349 2177 4401 2229
rect 4349 2113 4401 2165
rect 4349 2049 4401 2101
rect 4349 1985 4401 2037
rect 4349 1921 4401 1973
rect 4349 1857 4401 1909
rect 4349 1793 4401 1845
rect 4349 1729 4401 1781
rect 4349 1665 4401 1717
rect 4349 1601 4401 1653
rect 4349 1537 4401 1589
rect 4665 2177 4717 2229
rect 4665 2113 4717 2165
rect 4665 2049 4717 2101
rect 4665 1985 4717 2037
rect 4665 1921 4717 1973
rect 4665 1857 4717 1909
rect 4665 1793 4717 1845
rect 4665 1729 4717 1781
rect 4665 1665 4717 1717
rect 4665 1601 4717 1653
rect 4665 1537 4717 1589
rect 4981 2177 5033 2229
rect 4981 2113 5033 2165
rect 4981 2049 5033 2101
rect 4981 1985 5033 2037
rect 4981 1921 5033 1973
rect 4981 1857 5033 1909
rect 4981 1793 5033 1845
rect 4981 1729 5033 1781
rect 4981 1665 5033 1717
rect 4981 1601 5033 1653
rect 4981 1537 5033 1589
rect 5297 2177 5349 2229
rect 5297 2113 5349 2165
rect 5297 2049 5349 2101
rect 5297 1985 5349 2037
rect 5297 1921 5349 1973
rect 5297 1857 5349 1909
rect 5297 1793 5349 1845
rect 5297 1729 5349 1781
rect 5297 1665 5349 1717
rect 5297 1601 5349 1653
rect 5297 1537 5349 1589
rect 1663 338 1715 390
rect 1663 274 1715 326
rect 1663 210 1715 262
rect 1663 146 1715 198
rect 1663 82 1715 134
rect 1663 18 1715 70
rect 1663 -46 1715 6
rect 1663 -110 1715 -58
rect 1663 -174 1715 -122
rect 1663 -238 1715 -186
rect 1663 -302 1715 -250
rect 1979 338 2031 390
rect 1979 274 2031 326
rect 1979 210 2031 262
rect 1979 146 2031 198
rect 1979 82 2031 134
rect 1979 18 2031 70
rect 1979 -46 2031 6
rect 1979 -110 2031 -58
rect 1979 -174 2031 -122
rect 1979 -238 2031 -186
rect 1979 -302 2031 -250
rect 2295 338 2347 390
rect 2295 274 2347 326
rect 2295 210 2347 262
rect 2295 146 2347 198
rect 2295 82 2347 134
rect 2295 18 2347 70
rect 2295 -46 2347 6
rect 2295 -110 2347 -58
rect 2295 -174 2347 -122
rect 2295 -238 2347 -186
rect 2295 -302 2347 -250
rect 2611 338 2663 390
rect 2611 274 2663 326
rect 2611 210 2663 262
rect 2611 146 2663 198
rect 2611 82 2663 134
rect 2611 18 2663 70
rect 2611 -46 2663 6
rect 2611 -110 2663 -58
rect 2611 -174 2663 -122
rect 2611 -238 2663 -186
rect 2611 -302 2663 -250
rect 2927 338 2979 390
rect 2927 274 2979 326
rect 2927 210 2979 262
rect 2927 146 2979 198
rect 2927 82 2979 134
rect 2927 18 2979 70
rect 2927 -46 2979 6
rect 2927 -110 2979 -58
rect 2927 -174 2979 -122
rect 2927 -238 2979 -186
rect 2927 -302 2979 -250
rect 3243 338 3295 390
rect 3243 274 3295 326
rect 3243 210 3295 262
rect 3243 146 3295 198
rect 3243 82 3295 134
rect 3243 18 3295 70
rect 3243 -46 3295 6
rect 3243 -110 3295 -58
rect 3243 -174 3295 -122
rect 3243 -238 3295 -186
rect 3243 -302 3295 -250
rect 3559 338 3611 390
rect 3559 274 3611 326
rect 3559 210 3611 262
rect 3559 146 3611 198
rect 3559 82 3611 134
rect 3559 18 3611 70
rect 3559 -46 3611 6
rect 3559 -110 3611 -58
rect 3559 -174 3611 -122
rect 3559 -238 3611 -186
rect 3559 -302 3611 -250
rect 3875 338 3927 390
rect 3875 274 3927 326
rect 3875 210 3927 262
rect 3875 146 3927 198
rect 3875 82 3927 134
rect 3875 18 3927 70
rect 3875 -46 3927 6
rect 3875 -110 3927 -58
rect 3875 -174 3927 -122
rect 3875 -238 3927 -186
rect 3875 -302 3927 -250
rect 4191 338 4243 390
rect 4191 274 4243 326
rect 4191 210 4243 262
rect 4191 146 4243 198
rect 4191 82 4243 134
rect 4191 18 4243 70
rect 4191 -46 4243 6
rect 4191 -110 4243 -58
rect 4191 -174 4243 -122
rect 4191 -238 4243 -186
rect 4191 -302 4243 -250
rect 4507 338 4559 390
rect 4507 274 4559 326
rect 4507 210 4559 262
rect 4507 146 4559 198
rect 4507 82 4559 134
rect 4507 18 4559 70
rect 4507 -46 4559 6
rect 4507 -110 4559 -58
rect 4507 -174 4559 -122
rect 4507 -238 4559 -186
rect 4507 -302 4559 -250
rect 4823 338 4875 390
rect 4823 274 4875 326
rect 4823 210 4875 262
rect 4823 146 4875 198
rect 4823 82 4875 134
rect 4823 18 4875 70
rect 4823 -46 4875 6
rect 4823 -110 4875 -58
rect 4823 -174 4875 -122
rect 4823 -238 4875 -186
rect 4823 -302 4875 -250
rect 5139 338 5191 390
rect 5139 274 5191 326
rect 5139 210 5191 262
rect 5139 146 5191 198
rect 5139 82 5191 134
rect 5139 18 5191 70
rect 5139 -46 5191 6
rect 5139 -110 5191 -58
rect 5139 -174 5191 -122
rect 5139 -238 5191 -186
rect 5139 -302 5191 -250
rect 5455 338 5507 390
rect 5455 274 5507 326
rect 5455 210 5507 262
rect 5455 146 5507 198
rect 5455 82 5507 134
rect 5455 18 5507 70
rect 5455 -46 5507 6
rect 5455 -110 5507 -58
rect 5455 -174 5507 -122
rect 5455 -238 5507 -186
rect 5455 -302 5507 -250
rect 6081 2187 6261 2196
rect 6081 1577 6082 2187
rect 6082 1577 6260 2187
rect 6260 1577 6261 2187
rect 6081 1568 6261 1577
<< metal2 >>
rect 690 2229 6312 2260
rect 690 2185 1505 2229
rect 690 1557 744 2185
rect 924 2177 1505 2185
rect 1557 2177 1821 2229
rect 1873 2177 2137 2229
rect 2189 2177 2453 2229
rect 2505 2177 2769 2229
rect 2821 2177 3085 2229
rect 3137 2177 3401 2229
rect 3453 2177 3717 2229
rect 3769 2177 4033 2229
rect 4085 2177 4349 2229
rect 4401 2177 4665 2229
rect 4717 2177 4981 2229
rect 5033 2177 5297 2229
rect 5349 2196 6312 2229
rect 5349 2177 6081 2196
rect 924 2165 6081 2177
rect 924 2113 1505 2165
rect 1557 2113 1821 2165
rect 1873 2113 2137 2165
rect 2189 2113 2453 2165
rect 2505 2113 2769 2165
rect 2821 2113 3085 2165
rect 3137 2113 3401 2165
rect 3453 2113 3717 2165
rect 3769 2113 4033 2165
rect 4085 2113 4349 2165
rect 4401 2113 4665 2165
rect 4717 2113 4981 2165
rect 5033 2113 5297 2165
rect 5349 2113 6081 2165
rect 924 2101 6081 2113
rect 924 2049 1505 2101
rect 1557 2049 1821 2101
rect 1873 2049 2137 2101
rect 2189 2049 2453 2101
rect 2505 2049 2769 2101
rect 2821 2049 3085 2101
rect 3137 2049 3401 2101
rect 3453 2049 3717 2101
rect 3769 2049 4033 2101
rect 4085 2049 4349 2101
rect 4401 2049 4665 2101
rect 4717 2049 4981 2101
rect 5033 2049 5297 2101
rect 5349 2049 6081 2101
rect 924 2037 6081 2049
rect 924 1985 1505 2037
rect 1557 1985 1821 2037
rect 1873 1985 2137 2037
rect 2189 1985 2453 2037
rect 2505 1985 2769 2037
rect 2821 1985 3085 2037
rect 3137 1985 3401 2037
rect 3453 1985 3717 2037
rect 3769 1985 4033 2037
rect 4085 1985 4349 2037
rect 4401 1985 4665 2037
rect 4717 1985 4981 2037
rect 5033 1985 5297 2037
rect 5349 1985 6081 2037
rect 924 1973 6081 1985
rect 924 1921 1505 1973
rect 1557 1921 1821 1973
rect 1873 1921 2137 1973
rect 2189 1921 2453 1973
rect 2505 1921 2769 1973
rect 2821 1921 3085 1973
rect 3137 1921 3401 1973
rect 3453 1921 3717 1973
rect 3769 1921 4033 1973
rect 4085 1921 4349 1973
rect 4401 1921 4665 1973
rect 4717 1921 4981 1973
rect 5033 1921 5297 1973
rect 5349 1921 6081 1973
rect 924 1909 6081 1921
rect 924 1857 1505 1909
rect 1557 1857 1821 1909
rect 1873 1857 2137 1909
rect 2189 1857 2453 1909
rect 2505 1857 2769 1909
rect 2821 1857 3085 1909
rect 3137 1857 3401 1909
rect 3453 1857 3717 1909
rect 3769 1857 4033 1909
rect 4085 1857 4349 1909
rect 4401 1857 4665 1909
rect 4717 1857 4981 1909
rect 5033 1857 5297 1909
rect 5349 1857 6081 1909
rect 924 1845 6081 1857
rect 924 1793 1505 1845
rect 1557 1793 1821 1845
rect 1873 1793 2137 1845
rect 2189 1793 2453 1845
rect 2505 1793 2769 1845
rect 2821 1793 3085 1845
rect 3137 1793 3401 1845
rect 3453 1793 3717 1845
rect 3769 1793 4033 1845
rect 4085 1793 4349 1845
rect 4401 1793 4665 1845
rect 4717 1793 4981 1845
rect 5033 1793 5297 1845
rect 5349 1793 6081 1845
rect 924 1781 6081 1793
rect 924 1729 1505 1781
rect 1557 1729 1821 1781
rect 1873 1729 2137 1781
rect 2189 1729 2453 1781
rect 2505 1729 2769 1781
rect 2821 1729 3085 1781
rect 3137 1729 3401 1781
rect 3453 1729 3717 1781
rect 3769 1729 4033 1781
rect 4085 1729 4349 1781
rect 4401 1729 4665 1781
rect 4717 1729 4981 1781
rect 5033 1729 5297 1781
rect 5349 1729 6081 1781
rect 924 1717 6081 1729
rect 924 1665 1505 1717
rect 1557 1665 1821 1717
rect 1873 1665 2137 1717
rect 2189 1665 2453 1717
rect 2505 1665 2769 1717
rect 2821 1665 3085 1717
rect 3137 1665 3401 1717
rect 3453 1665 3717 1717
rect 3769 1665 4033 1717
rect 4085 1665 4349 1717
rect 4401 1665 4665 1717
rect 4717 1665 4981 1717
rect 5033 1665 5297 1717
rect 5349 1665 6081 1717
rect 924 1653 6081 1665
rect 924 1601 1505 1653
rect 1557 1601 1821 1653
rect 1873 1601 2137 1653
rect 2189 1601 2453 1653
rect 2505 1601 2769 1653
rect 2821 1601 3085 1653
rect 3137 1601 3401 1653
rect 3453 1601 3717 1653
rect 3769 1601 4033 1653
rect 4085 1601 4349 1653
rect 4401 1601 4665 1653
rect 4717 1601 4981 1653
rect 5033 1601 5297 1653
rect 5349 1601 6081 1653
rect 924 1589 6081 1601
rect 924 1557 1505 1589
rect 690 1537 1505 1557
rect 1557 1537 1821 1589
rect 1873 1537 2137 1589
rect 2189 1537 2453 1589
rect 2505 1537 2769 1589
rect 2821 1537 3085 1589
rect 3137 1537 3401 1589
rect 3453 1537 3717 1589
rect 3769 1537 4033 1589
rect 4085 1537 4349 1589
rect 4401 1537 4665 1589
rect 4717 1537 4981 1589
rect 5033 1537 5297 1589
rect 5349 1568 6081 1589
rect 6261 1568 6312 2196
rect 5349 1537 6312 1568
rect 690 1507 6312 1537
rect 1502 390 5510 424
rect 1502 338 1663 390
rect 1715 338 1979 390
rect 2031 338 2295 390
rect 2347 338 2611 390
rect 2663 338 2927 390
rect 2979 338 3243 390
rect 3295 338 3559 390
rect 3611 338 3875 390
rect 3927 338 4191 390
rect 4243 338 4507 390
rect 4559 338 4823 390
rect 4875 338 5139 390
rect 5191 338 5455 390
rect 5507 338 5510 390
rect 1502 326 5510 338
rect 1502 274 1663 326
rect 1715 274 1979 326
rect 2031 274 2295 326
rect 2347 274 2611 326
rect 2663 274 2927 326
rect 2979 274 3243 326
rect 3295 274 3559 326
rect 3611 274 3875 326
rect 3927 274 4191 326
rect 4243 274 4507 326
rect 4559 274 4823 326
rect 4875 274 5139 326
rect 5191 274 5455 326
rect 5507 274 5510 326
rect 1502 262 5510 274
rect 1502 210 1663 262
rect 1715 210 1979 262
rect 2031 210 2295 262
rect 2347 210 2611 262
rect 2663 210 2927 262
rect 2979 210 3243 262
rect 3295 210 3559 262
rect 3611 210 3875 262
rect 3927 210 4191 262
rect 4243 210 4507 262
rect 4559 210 4823 262
rect 4875 210 5139 262
rect 5191 210 5455 262
rect 5507 210 5510 262
rect 1502 198 5510 210
rect 1502 146 1663 198
rect 1715 146 1979 198
rect 2031 146 2295 198
rect 2347 146 2611 198
rect 2663 146 2927 198
rect 2979 146 3243 198
rect 3295 146 3559 198
rect 3611 146 3875 198
rect 3927 146 4191 198
rect 4243 146 4507 198
rect 4559 146 4823 198
rect 4875 146 5139 198
rect 5191 146 5455 198
rect 5507 146 5510 198
rect 1502 134 5510 146
rect 1502 82 1663 134
rect 1715 82 1979 134
rect 2031 82 2295 134
rect 2347 82 2611 134
rect 2663 82 2927 134
rect 2979 82 3243 134
rect 3295 82 3559 134
rect 3611 82 3875 134
rect 3927 82 4191 134
rect 4243 82 4507 134
rect 4559 82 4823 134
rect 4875 82 5139 134
rect 5191 82 5455 134
rect 5507 82 5510 134
rect 1502 70 5510 82
rect 1502 18 1663 70
rect 1715 18 1979 70
rect 2031 18 2295 70
rect 2347 18 2611 70
rect 2663 18 2927 70
rect 2979 18 3243 70
rect 3295 18 3559 70
rect 3611 18 3875 70
rect 3927 18 4191 70
rect 4243 18 4507 70
rect 4559 18 4823 70
rect 4875 18 5139 70
rect 5191 18 5455 70
rect 5507 18 5510 70
rect 1502 6 5510 18
rect 1502 -46 1663 6
rect 1715 -46 1979 6
rect 2031 -46 2295 6
rect 2347 -46 2611 6
rect 2663 -46 2927 6
rect 2979 -46 3243 6
rect 3295 -46 3559 6
rect 3611 -46 3875 6
rect 3927 -46 4191 6
rect 4243 -46 4507 6
rect 4559 -46 4823 6
rect 4875 -46 5139 6
rect 5191 -46 5455 6
rect 5507 -46 5510 6
rect 1502 -58 5510 -46
rect 1502 -110 1663 -58
rect 1715 -110 1979 -58
rect 2031 -110 2295 -58
rect 2347 -110 2611 -58
rect 2663 -110 2927 -58
rect 2979 -110 3243 -58
rect 3295 -110 3559 -58
rect 3611 -110 3875 -58
rect 3927 -110 4191 -58
rect 4243 -110 4507 -58
rect 4559 -110 4823 -58
rect 4875 -110 5139 -58
rect 5191 -110 5455 -58
rect 5507 -110 5510 -58
rect 1502 -122 5510 -110
rect 1502 -174 1663 -122
rect 1715 -174 1979 -122
rect 2031 -174 2295 -122
rect 2347 -174 2611 -122
rect 2663 -174 2927 -122
rect 2979 -174 3243 -122
rect 3295 -174 3559 -122
rect 3611 -174 3875 -122
rect 3927 -174 4191 -122
rect 4243 -174 4507 -122
rect 4559 -174 4823 -122
rect 4875 -174 5139 -122
rect 5191 -174 5455 -122
rect 5507 -174 5510 -122
rect 1502 -186 5510 -174
rect 1502 -238 1663 -186
rect 1715 -238 1979 -186
rect 2031 -238 2295 -186
rect 2347 -238 2611 -186
rect 2663 -238 2927 -186
rect 2979 -238 3243 -186
rect 3295 -238 3559 -186
rect 3611 -238 3875 -186
rect 3927 -238 4191 -186
rect 4243 -238 4507 -186
rect 4559 -238 4823 -186
rect 4875 -238 5139 -186
rect 5191 -238 5455 -186
rect 5507 -238 5510 -186
rect 1502 -250 5510 -238
rect 1502 -302 1663 -250
rect 1715 -302 1979 -250
rect 2031 -302 2295 -250
rect 2347 -302 2611 -250
rect 2663 -302 2927 -250
rect 2979 -302 3243 -250
rect 3295 -302 3559 -250
rect 3611 -302 3875 -250
rect 3927 -302 4191 -250
rect 4243 -302 4507 -250
rect 4559 -302 4823 -250
rect 4875 -302 5139 -250
rect 5191 -302 5455 -250
rect 5507 -302 5510 -250
rect 1502 -327 5510 -302
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_24
timestamp 1640969486
transform 1 0 1610 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_23
timestamp 1640969486
transform 1 0 1768 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_22
timestamp 1640969486
transform 1 0 1926 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_21
timestamp 1640969486
transform 1 0 2084 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_20
timestamp 1640969486
transform 1 0 2242 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_19
timestamp 1640969486
transform 1 0 2400 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_18
timestamp 1640969486
transform 1 0 2558 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_17
timestamp 1640969486
transform 1 0 2716 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_16
timestamp 1640969486
transform 1 0 2874 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_15
timestamp 1640969486
transform 1 0 3032 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_14
timestamp 1640969486
transform 1 0 3190 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_13
timestamp 1640969486
transform 1 0 3506 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_12
timestamp 1640969486
transform 1 0 3348 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_11
timestamp 1640969486
transform 1 0 3822 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_10
timestamp 1640969486
transform 1 0 3664 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_9
timestamp 1640969486
transform 1 0 4138 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_8
timestamp 1640969486
transform 1 0 3980 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_7
timestamp 1640969486
transform 1 0 4454 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_6
timestamp 1640969486
transform 1 0 4296 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_5
timestamp 1640969486
transform 1 0 4770 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_4
timestamp 1640969486
transform 1 0 4612 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_3
timestamp 1640969486
transform 1 0 4928 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_2
timestamp 1640969486
transform 1 0 5086 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_1
timestamp 1640969486
transform 1 0 5244 0 1 870
box -144 -1482 144 1482
use sky130_fd_pr__pfet_01v8_lvt_WFBLZ7  sky130_fd_pr__pfet_01v8_lvt_WFBLZ7_0
timestamp 1640969486
transform 1 0 5402 0 1 870
box -144 -1482 144 1482
<< labels >>
flabel metal2 s 1048 1826 1048 1826 0 FreeSans 2000 0 0 0 S
port 1 nsew
flabel metal2 s 1614 -57 1614 -57 0 FreeSans 2000 0 0 0 D
port 2 nsew
flabel metal1 s 1334 544 1334 544 0 FreeSans 2000 0 0 0 G
port 3 nsew
<< end >>
