magic
tech sky130A
magscale 1 2
timestamp 1640969486
<< nwell >>
rect -774 -1381 23357 1700
rect -774 -1702 24510 -1381
rect -774 -1789 5028 -1702
rect 7430 -1789 24510 -1702
rect 12870 -2502 24510 -1789
rect 12870 -3140 12888 -2502
rect 13002 -2696 13150 -2502
rect 18686 -2728 18830 -2502
<< pwell >>
rect -134 -3052 110 -2176
rect 6054 -3366 6288 -2396
<< psubdiff >>
rect -108 -2256 84 -2202
rect -108 -2970 -64 -2256
rect 38 -2970 84 -2256
rect -108 -3026 84 -2970
rect 6080 -2487 6262 -2422
rect 6080 -3269 6117 -2487
rect 6219 -3269 6262 -2487
rect 6080 -3340 6262 -3269
<< mvnsubdiff >>
rect -66 1039 222 1212
rect -66 325 -12 1039
rect 158 501 222 1039
rect 5694 676 5804 720
rect 5694 642 5727 676
rect 5761 642 5804 676
rect 5694 608 5804 642
rect 5694 574 5727 608
rect 5761 574 5804 608
rect 5694 540 5804 574
rect 5694 506 5727 540
rect 5761 506 5804 540
rect 158 325 228 501
rect -66 277 228 325
rect -58 198 228 277
rect 5694 472 5804 506
rect 5694 438 5727 472
rect 5761 438 5804 472
rect 5694 404 5804 438
rect 5694 370 5727 404
rect 5761 370 5804 404
rect 5694 336 5804 370
rect 5694 302 5727 336
rect 5761 302 5804 336
rect 5694 248 5804 302
rect 11286 716 11444 764
rect 11286 682 11345 716
rect 11379 682 11444 716
rect 11286 648 11444 682
rect 11286 614 11345 648
rect 11379 614 11444 648
rect 11286 580 11444 614
rect 11286 546 11345 580
rect 11379 546 11444 580
rect 11286 512 11444 546
rect 11286 478 11345 512
rect 11379 478 11444 512
rect 11286 444 11444 478
rect 11286 410 11345 444
rect 11379 410 11444 444
rect 11286 376 11444 410
rect 11286 342 11345 376
rect 11379 342 11444 376
rect 11286 308 11444 342
rect 11286 274 11345 308
rect 11379 274 11444 308
rect 11286 230 11444 274
rect -58 -44 2009 198
rect -8 -47 2009 -44
rect -232 -688 -70 -618
rect -232 -1198 -206 -688
rect -104 -1198 -70 -688
rect -232 -1276 -70 -1198
rect 5494 -817 5606 -784
rect 5494 -851 5528 -817
rect 5562 -851 5606 -817
rect 5494 -885 5606 -851
rect 5494 -919 5528 -885
rect 5562 -919 5606 -885
rect 5494 -953 5606 -919
rect 5494 -987 5528 -953
rect 5562 -987 5606 -953
rect 5494 -1021 5606 -987
rect 5494 -1055 5528 -1021
rect 5562 -1055 5606 -1021
rect 5494 -1089 5606 -1055
rect 5494 -1123 5528 -1089
rect 5562 -1123 5606 -1089
rect 5494 -1157 5606 -1123
rect 5494 -1191 5528 -1157
rect 5562 -1191 5606 -1157
rect 5494 -1220 5606 -1191
rect 16774 -837 16872 -770
rect 16774 -871 16803 -837
rect 16837 -871 16872 -837
rect 16774 -905 16872 -871
rect 16774 -939 16803 -905
rect 16837 -939 16872 -905
rect 16774 -973 16872 -939
rect 16774 -1007 16803 -973
rect 16837 -1007 16872 -973
rect 16774 -1041 16872 -1007
rect 16774 -1075 16803 -1041
rect 16837 -1075 16872 -1041
rect 16774 -1109 16872 -1075
rect 16774 -1143 16803 -1109
rect 16837 -1143 16872 -1109
rect 16774 -1202 16872 -1143
rect 22422 -790 22546 -744
rect 22422 -824 22468 -790
rect 22502 -824 22546 -790
rect 22422 -858 22546 -824
rect 22422 -892 22468 -858
rect 22502 -892 22546 -858
rect 22422 -926 22546 -892
rect 22422 -960 22468 -926
rect 22502 -960 22546 -926
rect 22422 -994 22546 -960
rect 22422 -1028 22468 -994
rect 22502 -1028 22546 -994
rect 22422 -1062 22546 -1028
rect 22422 -1096 22468 -1062
rect 22502 -1096 22546 -1062
rect 22422 -1130 22546 -1096
rect 22422 -1164 22468 -1130
rect 22502 -1164 22546 -1130
rect 22422 -1198 22546 -1164
rect 22422 -1232 22468 -1198
rect 22502 -1232 22546 -1198
rect 22422 -1306 22546 -1232
rect 13002 -2347 13150 -2302
rect 13002 -2381 13059 -2347
rect 13093 -2381 13150 -2347
rect 13002 -2415 13150 -2381
rect 13002 -2449 13059 -2415
rect 13093 -2449 13150 -2415
rect 13002 -2483 13150 -2449
rect 13002 -2517 13059 -2483
rect 13093 -2517 13150 -2483
rect 13002 -2551 13150 -2517
rect 13002 -2585 13059 -2551
rect 13093 -2585 13150 -2551
rect 13002 -2619 13150 -2585
rect 13002 -2653 13059 -2619
rect 13093 -2653 13150 -2619
rect 13002 -2696 13150 -2653
rect 18702 -2369 18804 -2330
rect 18702 -2403 18734 -2369
rect 18768 -2403 18804 -2369
rect 18702 -2437 18804 -2403
rect 18702 -2471 18734 -2437
rect 18768 -2471 18804 -2437
rect 18702 -2505 18804 -2471
rect 18702 -2539 18734 -2505
rect 18768 -2539 18804 -2505
rect 18702 -2573 18804 -2539
rect 18702 -2607 18734 -2573
rect 18768 -2607 18804 -2573
rect 18702 -2641 18804 -2607
rect 18702 -2675 18734 -2641
rect 18768 -2675 18804 -2641
rect 18702 -2704 18804 -2675
<< psubdiffcont >>
rect -64 -2970 38 -2256
rect 6117 -3269 6219 -2487
<< mvnsubdiffcont >>
rect -12 325 158 1039
rect 5727 642 5761 676
rect 5727 574 5761 608
rect 5727 506 5761 540
rect 5727 438 5761 472
rect 5727 370 5761 404
rect 5727 302 5761 336
rect 11345 682 11379 716
rect 11345 614 11379 648
rect 11345 546 11379 580
rect 11345 478 11379 512
rect 11345 410 11379 444
rect 11345 342 11379 376
rect 11345 274 11379 308
rect -206 -1198 -104 -688
rect 5528 -851 5562 -817
rect 5528 -919 5562 -885
rect 5528 -987 5562 -953
rect 5528 -1055 5562 -1021
rect 5528 -1123 5562 -1089
rect 5528 -1191 5562 -1157
rect 16803 -871 16837 -837
rect 16803 -939 16837 -905
rect 16803 -1007 16837 -973
rect 16803 -1075 16837 -1041
rect 16803 -1143 16837 -1109
rect 22468 -824 22502 -790
rect 22468 -892 22502 -858
rect 22468 -960 22502 -926
rect 22468 -1028 22502 -994
rect 22468 -1096 22502 -1062
rect 22468 -1164 22502 -1130
rect 22468 -1232 22502 -1198
rect 13059 -2381 13093 -2347
rect 13059 -2449 13093 -2415
rect 13059 -2517 13093 -2483
rect 13059 -2585 13093 -2551
rect 13059 -2653 13093 -2619
rect 18734 -2403 18768 -2369
rect 18734 -2471 18768 -2437
rect 18734 -2539 18768 -2505
rect 18734 -2607 18768 -2573
rect 18734 -2675 18768 -2641
<< locali >>
rect -58 1504 21652 2590
rect -58 1494 22678 1504
rect -58 1218 22682 1494
rect -58 1212 21652 1218
rect -66 1210 21652 1212
rect -66 1039 222 1210
rect -66 486 -12 1039
rect -278 325 -12 486
rect 158 501 222 1039
rect 5688 676 5816 1210
rect 5688 642 5727 676
rect 5761 642 5816 676
rect 5688 608 5816 642
rect 5688 574 5727 608
rect 5761 574 5816 608
rect 5688 540 5816 574
rect 5688 506 5727 540
rect 5761 506 5816 540
rect 158 325 228 501
rect -278 198 228 325
rect 5688 472 5816 506
rect 5688 438 5727 472
rect 5761 438 5816 472
rect 5688 404 5816 438
rect 5688 370 5727 404
rect 5761 370 5816 404
rect 5688 336 5816 370
rect 5688 302 5727 336
rect 5761 302 5816 336
rect -278 -47 2009 198
rect 5688 196 5816 302
rect 11238 716 11498 1210
rect 11238 682 11345 716
rect 11379 682 11498 716
rect 11238 648 11498 682
rect 11238 614 11345 648
rect 11379 614 11498 648
rect 11238 580 11498 614
rect 11238 546 11345 580
rect 11379 546 11498 580
rect 11238 512 11498 546
rect 11238 478 11345 512
rect 11379 478 11498 512
rect 11238 444 11498 478
rect 11238 410 11345 444
rect 11379 410 11498 444
rect 11238 376 11498 410
rect 11238 342 11345 376
rect 11379 342 11498 376
rect 11238 308 11498 342
rect 11238 274 11345 308
rect 11379 274 11498 308
rect 11238 216 11498 274
rect -278 -638 20 -47
rect 4769 -49 6437 196
rect 9383 2 13146 216
rect 16950 211 17210 1210
rect 16046 -85 17210 211
rect 16950 -100 17210 -85
rect -272 -688 -30 -638
rect -272 -1198 -206 -688
rect -104 -1198 -30 -688
rect -272 -1326 -30 -1198
rect 5474 -817 5626 -750
rect 5474 -851 5528 -817
rect 5562 -851 5626 -817
rect 5474 -885 5626 -851
rect 5474 -919 5528 -885
rect 5562 -919 5626 -885
rect 5474 -953 5626 -919
rect 5474 -987 5528 -953
rect 5562 -987 5626 -953
rect 5474 -1021 5626 -987
rect 5474 -1055 5528 -1021
rect 5562 -1055 5626 -1021
rect 5474 -1089 5626 -1055
rect 5474 -1123 5528 -1089
rect 5562 -1123 5626 -1089
rect 5474 -1157 5626 -1123
rect 5474 -1191 5528 -1157
rect 5562 -1191 5626 -1157
rect 5474 -1248 5626 -1191
rect 16746 -837 16900 -746
rect 22394 -790 22682 1218
rect 22394 -816 22468 -790
rect 16746 -871 16803 -837
rect 16837 -871 16900 -837
rect 16746 -905 16900 -871
rect 16746 -939 16803 -905
rect 16837 -939 16900 -905
rect 16746 -973 16900 -939
rect 16746 -1007 16803 -973
rect 16837 -1007 16900 -973
rect 16746 -1041 16900 -1007
rect 16746 -1075 16803 -1041
rect 16837 -1075 16900 -1041
rect 16746 -1109 16900 -1075
rect 16746 -1143 16803 -1109
rect 16837 -1143 16900 -1109
rect 16746 -1234 16900 -1143
rect 22406 -824 22468 -816
rect 22502 -816 22682 -790
rect 22502 -824 22566 -816
rect 22406 -858 22566 -824
rect 22406 -892 22468 -858
rect 22502 -892 22566 -858
rect 22406 -926 22566 -892
rect 22406 -960 22468 -926
rect 22502 -960 22566 -926
rect 22406 -994 22566 -960
rect 22406 -1028 22468 -994
rect 22502 -1028 22566 -994
rect 22406 -1062 22566 -1028
rect 22406 -1096 22468 -1062
rect 22502 -1096 22566 -1062
rect 22406 -1130 22566 -1096
rect 22406 -1164 22468 -1130
rect 22502 -1164 22566 -1130
rect 22406 -1198 22566 -1164
rect 22406 -1232 22468 -1198
rect 22502 -1232 22566 -1198
rect 22406 -1338 22566 -1232
rect -146 -2256 130 -2158
rect -146 -2970 -64 -2256
rect 38 -2970 130 -2256
rect 13002 -2347 13150 -2302
rect -146 -2974 130 -2970
rect 6046 -2487 6296 -2366
rect -186 -3824 178 -2974
rect 6046 -3269 6117 -2487
rect 6219 -3269 6296 -2487
rect 13002 -2381 13059 -2347
rect 13093 -2381 13150 -2347
rect 13002 -2415 13150 -2381
rect 13002 -2449 13059 -2415
rect 13093 -2449 13150 -2415
rect 13002 -2483 13150 -2449
rect 13002 -2517 13059 -2483
rect 13093 -2517 13150 -2483
rect 13002 -2551 13150 -2517
rect 13002 -2585 13059 -2551
rect 13093 -2585 13150 -2551
rect 13002 -2619 13150 -2585
rect 13002 -2653 13059 -2619
rect 13093 -2653 13150 -2619
rect 13002 -2696 13150 -2653
rect 18686 -2369 18830 -2310
rect 18686 -2403 18734 -2369
rect 18768 -2403 18830 -2369
rect 18686 -2437 18830 -2403
rect 18686 -2471 18734 -2437
rect 18768 -2471 18830 -2437
rect 18686 -2505 18830 -2471
rect 18686 -2539 18734 -2505
rect 18768 -2539 18830 -2505
rect 18686 -2573 18830 -2539
rect 18686 -2607 18734 -2573
rect 18768 -2607 18830 -2573
rect 18686 -2641 18830 -2607
rect 18686 -2675 18734 -2641
rect 18768 -2675 18830 -2641
rect 18686 -2728 18830 -2675
rect 6046 -3374 6296 -3269
rect -186 -4048 966 -3824
rect 10602 -3920 10866 -2850
rect 10602 -4098 10641 -3920
rect 10819 -4098 10866 -3920
rect 10602 -4166 10866 -4098
rect 9524 -5006 10072 -4710
rect 12164 -5006 12640 -2934
rect 13334 -5006 14586 -4540
rect 15374 -5006 15692 -4276
rect -142 -5780 19804 -5006
<< viali >>
rect 10641 -4098 10819 -3920
<< metal1 >>
rect 15408 1072 15844 1092
rect 15400 1027 15844 1072
rect 3161 990 8624 991
rect 3161 787 14289 990
rect 3161 781 8624 787
rect 15400 783 15447 1027
rect 15755 783 15844 1027
rect 15400 722 15844 783
rect 15400 694 15826 722
rect 6645 664 7397 692
rect 2192 571 2755 625
rect 2192 391 2237 571
rect 2673 391 2755 571
rect 2192 325 2755 391
rect 6645 356 6718 664
rect 7282 356 7397 664
rect 6645 331 7397 356
rect 13302 -159 14564 -78
rect 8246 -581 8734 -546
rect 8246 -697 8293 -581
rect 8665 -697 8734 -581
rect 8246 -732 8734 -697
rect 13302 -659 13391 -159
rect 14467 -659 14564 -159
rect 15736 -204 15952 582
rect 15736 -259 17870 -204
rect 15736 -370 17439 -259
rect 15742 -439 17439 -370
rect 17811 -439 17870 -259
rect 15742 -512 17870 -439
rect 12064 -766 12726 -712
rect 13302 -714 14564 -659
rect 1825 -943 2590 -923
rect 1825 -1123 1898 -943
rect 2462 -1123 2590 -943
rect 12064 -1074 12131 -766
rect 12695 -1074 12726 -766
rect 12064 -1092 12726 -1074
rect 15412 -801 15798 -758
rect 15412 -1045 15486 -801
rect 15730 -1045 15798 -801
rect 15412 -1092 15798 -1045
rect 1825 -1155 2590 -1123
rect 1358 -2753 1812 -2712
rect 1358 -2933 1391 -2753
rect 1763 -2933 1812 -2753
rect 2258 -2806 2872 -1258
rect 5028 -1776 7430 -1702
rect 5028 -2214 7442 -1776
rect 5046 -2566 5620 -2214
rect 6868 -2548 7442 -2214
rect 11806 -2498 12048 -1244
rect 13768 -1911 14918 -1814
rect 13768 -2155 13810 -1911
rect 14822 -2155 14918 -1911
rect 13768 -2202 14918 -2155
rect 17392 -2406 17862 -2338
rect 3368 -2708 4086 -2676
rect 1358 -2976 1812 -2933
rect 3368 -2888 3419 -2708
rect 3983 -2888 4086 -2708
rect 3368 -2944 4086 -2888
rect 8304 -2684 8742 -2652
rect 8304 -2864 8388 -2684
rect 8696 -2864 8742 -2684
rect 11812 -2696 12038 -2498
rect 17392 -2586 17477 -2406
rect 17785 -2586 17862 -2406
rect 17392 -2642 17862 -2586
rect 8304 -2926 8742 -2864
rect 11712 -2798 12038 -2696
rect 11712 -2972 12030 -2798
rect 18784 -3364 19198 -2960
rect 18770 -3706 22220 -3364
rect 10544 -3920 10938 -3820
rect 10544 -4098 10641 -3920
rect 10819 -4098 10938 -3920
rect 210 -4220 880 -4130
rect 210 -4720 267 -4220
rect 767 -4720 880 -4220
rect 10544 -4488 10938 -4098
rect 14042 -4228 15334 -4056
rect 18784 -4236 19198 -3706
rect 8068 -4670 9660 -4494
rect 10216 -4658 10942 -4488
rect 210 -4780 880 -4720
<< via1 >>
rect 15447 783 15755 1027
rect 2237 391 2673 571
rect 6718 356 7282 664
rect 8293 -697 8665 -581
rect 13391 -659 14467 -159
rect 17439 -439 17811 -259
rect 1898 -1123 2462 -943
rect 12131 -1074 12695 -766
rect 15486 -1045 15730 -801
rect 1391 -2933 1763 -2753
rect 13810 -2155 14822 -1911
rect 3419 -2888 3983 -2708
rect 8388 -2864 8696 -2684
rect 17477 -2586 17785 -2406
rect 267 -4720 767 -4220
<< metal2 >>
rect 15380 1027 15876 1118
rect 15380 783 15447 1027
rect 15755 783 15876 1027
rect 6584 664 7477 753
rect 1849 571 2798 637
rect 1849 391 2237 571
rect 2673 391 2798 571
rect 1849 288 2798 391
rect 6584 356 6718 664
rect 7282 356 7477 664
rect 1849 -892 2541 288
rect 6584 282 7477 356
rect 6665 -94 7396 282
rect 6665 -444 12808 -94
rect 13276 -159 14676 -18
rect 6665 -462 7396 -444
rect 8136 -538 8800 -506
rect 8136 -754 8210 -538
rect 8746 -754 8800 -538
rect 8136 -794 8800 -754
rect 12002 -766 12799 -444
rect 1770 -943 2632 -892
rect 1770 -1123 1898 -943
rect 2462 -1123 2632 -943
rect 12002 -1074 12131 -766
rect 12695 -1074 12799 -766
rect 12002 -1104 12799 -1074
rect 13276 -659 13391 -159
rect 14467 -659 14676 -159
rect 1770 -1198 2632 -1123
rect 13276 -1578 14676 -659
rect 15380 -801 15876 783
rect 15380 -1045 15486 -801
rect 15730 -1045 15876 -801
rect 15380 -1142 15876 -1045
rect 17346 -259 17932 -178
rect 17346 -439 17439 -259
rect 17811 -439 17932 -259
rect 4066 -1586 14676 -1578
rect 3340 -1688 14676 -1586
rect 3340 -1911 15002 -1688
rect 3340 -2155 13810 -1911
rect 14822 -2155 15002 -1911
rect 3340 -2220 15002 -2155
rect 3340 -2224 14652 -2220
rect 1306 -2753 1840 -2694
rect 1306 -2933 1391 -2753
rect 1763 -2933 1840 -2753
rect 3340 -2708 4186 -2224
rect 17346 -2406 17932 -439
rect 17346 -2586 17477 -2406
rect 17785 -2586 17932 -2406
rect 3340 -2824 3419 -2708
rect 1306 -4086 1840 -2933
rect 3348 -2888 3419 -2824
rect 3983 -2824 4186 -2708
rect 8172 -2649 8774 -2648
rect 3983 -2888 4184 -2824
rect 3348 -2958 4184 -2888
rect 8172 -2865 8348 -2649
rect 8724 -2865 8774 -2649
rect 17346 -2672 17932 -2586
rect 8172 -2966 8774 -2865
rect 180 -4220 1840 -4086
rect 180 -4720 267 -4220
rect 767 -4720 1840 -4220
rect 180 -4828 1840 -4720
<< via2 >>
rect 8210 -581 8746 -538
rect 8210 -697 8293 -581
rect 8293 -697 8665 -581
rect 8665 -697 8746 -581
rect 8210 -754 8746 -697
rect 8348 -2684 8724 -2649
rect 8348 -2864 8388 -2684
rect 8388 -2864 8696 -2684
rect 8696 -2864 8724 -2684
rect 8348 -2865 8724 -2864
<< metal3 >>
rect 8088 -538 8830 -488
rect 8088 -754 8210 -538
rect 8746 -754 8830 -538
rect 8088 -2649 8830 -754
rect 8088 -2832 8348 -2649
rect 8090 -2865 8348 -2832
rect 8724 -2832 8830 -2649
rect 8724 -2865 8824 -2832
rect 8090 -2994 8824 -2865
use sky130_fd_pr__res_xhigh_po_0p35_6WVZEH  sky130_fd_pr__res_xhigh_po_0p35_6WVZEH_0
timestamp 1640969486
transform 0 -1 9788 1 0 -4584
box -191 -723 191 723
use BJT  BJT_0
timestamp 1640969486
transform 1 0 2162 0 1 -3784
box 0 -1342 6708 -2
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1640969486
transform 1 0 -160 0 1 -5138
box 0 0 1340 1340
use sky130_fd_pr__res_xhigh_po_0p35_47C2TB  sky130_fd_pr__res_xhigh_po_0p35_47C2TB_0
timestamp 1640969486
transform 0 -1 17079 1 0 -4156
box -191 -2268 191 2268
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0
timestamp 1640969486
transform 1 0 13304 0 1 -4796
box 0 0 1340 1340
use bgr_nmos  bgr_nmos_1
timestamp 1640969486
transform -1 0 11819 0 1 -3058
box -28 -123 5372 578
use bgr_nmos  bgr_nmos_0
timestamp 1640969486
transform 1 0 515 0 1 -3058
box -28 -123 5372 578
use bgr_pmos2  bgr_pmos2_2
timestamp 1640969486
transform 1 0 16209 0 1 -2598
box -3323 -542 8317 579
use bgr_pmos2  bgr_pmos2_0
timestamp 1640969486
transform -1 0 19374 0 1 -1091
box -3323 -542 8317 579
use bgr_pmos2  bgr_pmos2_1
timestamp 1640969486
transform 1 0 2997 0 1 -1091
box -3323 -542 8317 579
use bgr_pmos  bgr_pmos_0
timestamp 1640969486
transform -1 0 13932 0 1 380
box -3322 -380 2686 564
use bgr_pmos  bgr_pmos_1
timestamp 1640969486
transform 1 0 8815 0 1 380
box -3322 -380 2686 564
use bgr_pmos  bgr_pmos_2
timestamp 1640969486
transform -1 0 2686 0 1 380
box -3322 -380 2686 564
<< labels >>
flabel locali s 4296 -5516 4296 -5516 0 FreeSans 2500 0 0 0 VSS
port 1 nsew
flabel locali s 6538 1978 6538 1978 0 FreeSans 2500 0 0 0 VDD
port 2 nsew
flabel metal1 s 21846 -3476 21846 -3476 0 FreeSans 2500 0 0 0 VREF
port 3 nsew
<< end >>
