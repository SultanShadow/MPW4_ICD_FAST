magic
tech sky130A
magscale 1 2
timestamp 1640969486
<< nwell >>
rect 3788 2096 3822 2876
rect 14120 2390 14154 2930
rect 3872 2262 3922 2312
<< pwell >>
rect 4746 1490 4832 1710
rect 9060 1478 9146 1698
rect 9780 1470 9866 1690
rect 14094 1458 14180 1678
<< psubdiff >>
rect 4772 1516 4806 1684
rect 9086 1504 9120 1672
rect 9806 1496 9840 1664
rect 14120 1484 14154 1652
<< nsubdiff >>
rect 3788 2096 3822 2876
rect 14120 2390 14154 2930
<< poly >>
rect 3872 2262 3922 2312
rect 4852 1788 4912 1860
rect 8968 1786 9028 1858
rect 9880 1778 9952 1862
rect 4854 1334 4914 1406
rect 8970 1334 9030 1406
<< locali >>
rect 3788 2136 3822 2876
rect 4034 2794 4282 2938
rect 4088 2334 4336 2478
rect 14120 2390 14154 2930
rect 3788 2133 3858 2136
rect 3788 2099 3810 2133
rect 3844 2099 3858 2133
rect 3788 2096 3858 2099
rect 9180 2117 9744 2120
rect 9180 2083 9193 2117
rect 9227 2083 9265 2117
rect 9299 2083 9337 2117
rect 9371 2083 9409 2117
rect 9443 2083 9481 2117
rect 9515 2083 9553 2117
rect 9587 2083 9625 2117
rect 9659 2083 9697 2117
rect 9731 2083 9744 2117
rect 9180 2080 9744 2083
rect 9086 1926 9840 2018
rect 4772 1516 4806 1684
rect 9086 1504 9120 1672
rect 9806 1496 9840 1664
rect 11718 1636 12618 1772
rect 14120 1484 14154 1652
rect 5416 736 6316 872
rect 8978 680 9024 694
rect 3794 618 3812 652
rect 3846 618 3864 652
rect 8978 646 8984 680
rect 9018 646 9024 680
rect 8978 632 9024 646
<< viali >>
rect 3810 2099 3844 2133
rect 9193 2083 9227 2117
rect 9265 2083 9299 2117
rect 9337 2083 9371 2117
rect 9409 2083 9443 2117
rect 9481 2083 9515 2117
rect 9553 2083 9587 2117
rect 9625 2083 9659 2117
rect 9697 2083 9731 2117
rect 3812 618 3846 652
rect 8984 646 9018 680
<< metal1 >>
rect 3850 2769 3934 2794
rect 3850 2717 3872 2769
rect 3924 2717 3934 2769
rect 3850 2692 3934 2717
rect 14008 2714 14062 2778
rect 5100 2684 5812 2688
rect 5100 2632 5108 2684
rect 5160 2632 5172 2684
rect 5224 2632 5236 2684
rect 5288 2632 5300 2684
rect 5352 2632 5364 2684
rect 5416 2632 5428 2684
rect 5480 2632 5492 2684
rect 5544 2632 5556 2684
rect 5608 2632 5620 2684
rect 5672 2632 5684 2684
rect 5736 2632 5748 2684
rect 5800 2632 5812 2684
rect 5100 2608 5812 2632
rect 3862 2314 3932 2328
rect 3862 2262 3874 2314
rect 3926 2262 3932 2314
rect 3862 2252 3932 2262
rect 14010 2254 14064 2318
rect 7234 2226 7946 2230
rect 3792 2158 3886 2178
rect 3790 2133 3886 2158
rect 3790 2099 3810 2133
rect 3844 2099 3886 2133
rect 7234 2174 7275 2226
rect 7327 2174 7339 2226
rect 7391 2174 7403 2226
rect 7455 2174 7467 2226
rect 7519 2174 7531 2226
rect 7583 2174 7595 2226
rect 7647 2174 7659 2226
rect 7711 2174 7723 2226
rect 7775 2174 7787 2226
rect 7839 2174 7851 2226
rect 7903 2174 7946 2226
rect 7234 2128 7946 2174
rect 3790 1862 3886 2099
rect 9164 2117 9760 2126
rect 9164 2083 9193 2117
rect 9227 2083 9265 2117
rect 9299 2083 9337 2117
rect 9371 2083 9409 2117
rect 9443 2083 9481 2117
rect 9515 2083 9553 2117
rect 9587 2083 9625 2117
rect 9659 2083 9697 2117
rect 9731 2083 9760 2117
rect 5094 1930 5816 1950
rect 5094 1878 5109 1930
rect 5161 1878 5173 1930
rect 5225 1878 5237 1930
rect 5289 1878 5301 1930
rect 5353 1878 5365 1930
rect 5417 1878 5429 1930
rect 5481 1878 5493 1930
rect 5545 1878 5557 1930
rect 5609 1878 5621 1930
rect 5673 1878 5685 1930
rect 5737 1878 5749 1930
rect 5801 1878 5816 1930
rect 5094 1870 5816 1878
rect 9164 1862 9760 2083
rect 10630 1883 11404 1888
rect 10630 1882 10639 1883
rect 3790 1860 4908 1862
rect 3790 1788 4912 1860
rect 3790 1786 4908 1788
rect 3790 964 3886 1786
rect 8974 1784 9950 1862
rect 10614 1831 10639 1882
rect 10691 1831 10703 1883
rect 10755 1831 10767 1883
rect 10819 1831 10831 1883
rect 10883 1831 10895 1883
rect 10947 1831 10959 1883
rect 11011 1831 11023 1883
rect 11075 1831 11087 1883
rect 11139 1831 11151 1883
rect 11203 1831 11215 1883
rect 11267 1831 11279 1883
rect 11331 1831 11343 1883
rect 11395 1882 11404 1883
rect 11395 1831 11426 1882
rect 10614 1820 11426 1831
rect 14010 1794 14064 1858
rect 9164 1782 9760 1784
rect 6080 1772 6130 1774
rect 5182 1747 6130 1772
rect 5182 1695 5204 1747
rect 5256 1695 5268 1747
rect 5320 1695 5332 1747
rect 5384 1695 5396 1747
rect 5448 1695 5460 1747
rect 5512 1695 5524 1747
rect 5576 1695 5588 1747
rect 5640 1695 5652 1747
rect 5704 1695 5716 1747
rect 5768 1695 5780 1747
rect 5832 1695 5844 1747
rect 5896 1695 5908 1747
rect 5960 1695 5972 1747
rect 6024 1695 6036 1747
rect 6088 1695 6130 1747
rect 5182 1654 6130 1695
rect 5182 1648 6102 1654
rect 5152 1491 6136 1522
rect 5152 1439 5168 1491
rect 5220 1439 5232 1491
rect 5284 1439 5296 1491
rect 5348 1439 5360 1491
rect 5412 1439 5424 1491
rect 5476 1439 5488 1491
rect 5540 1439 5552 1491
rect 5604 1439 5616 1491
rect 5668 1439 5680 1491
rect 5732 1439 5744 1491
rect 5796 1439 5808 1491
rect 5860 1439 5872 1491
rect 5924 1439 5936 1491
rect 5988 1439 6000 1491
rect 6052 1439 6064 1491
rect 6116 1439 6136 1491
rect 5152 1424 6136 1439
rect 10602 1484 11454 1502
rect 6338 1436 6928 1438
rect 5164 1418 6120 1424
rect 4854 1334 4914 1406
rect 6338 1384 6391 1436
rect 6443 1384 6455 1436
rect 6507 1384 6519 1436
rect 6571 1384 6583 1436
rect 6635 1384 6647 1436
rect 6699 1384 6711 1436
rect 6763 1384 6775 1436
rect 6827 1384 6839 1436
rect 6891 1384 6928 1436
rect 10602 1432 10644 1484
rect 10696 1432 10708 1484
rect 10760 1432 10772 1484
rect 10824 1432 10836 1484
rect 10888 1432 10900 1484
rect 10952 1432 10964 1484
rect 11016 1432 11028 1484
rect 11080 1432 11092 1484
rect 11144 1432 11156 1484
rect 11208 1432 11220 1484
rect 11272 1432 11284 1484
rect 11336 1432 11348 1484
rect 11400 1432 11454 1484
rect 10616 1428 11428 1432
rect 6338 1372 6928 1384
rect 8974 1394 9950 1404
rect 7222 1356 7978 1378
rect 4028 1304 4294 1330
rect 7222 1304 7256 1356
rect 7308 1304 7320 1356
rect 7372 1304 7384 1356
rect 7436 1304 7448 1356
rect 7500 1304 7512 1356
rect 7564 1304 7576 1356
rect 7628 1304 7640 1356
rect 7692 1304 7704 1356
rect 7756 1304 7768 1356
rect 7820 1304 7832 1356
rect 7884 1304 7896 1356
rect 7948 1304 7978 1356
rect 8974 1342 9236 1394
rect 9288 1342 9300 1394
rect 9352 1342 9364 1394
rect 9416 1342 9428 1394
rect 9480 1342 9492 1394
rect 9544 1342 9556 1394
rect 9608 1342 9620 1394
rect 9672 1342 9950 1394
rect 8974 1334 9950 1342
rect 14010 1332 14064 1396
rect 4028 1291 5162 1304
rect 7222 1296 7978 1304
rect 11712 1297 12594 1304
rect 4028 1239 4060 1291
rect 4112 1239 4124 1291
rect 4176 1239 4188 1291
rect 4240 1239 5162 1291
rect 11712 1282 11743 1297
rect 4028 1212 5162 1239
rect 11690 1245 11743 1282
rect 11795 1245 11807 1297
rect 11859 1245 11871 1297
rect 11923 1245 11935 1297
rect 11987 1245 11999 1297
rect 12051 1245 12063 1297
rect 12115 1245 12127 1297
rect 12179 1245 12191 1297
rect 12243 1245 12255 1297
rect 12307 1245 12319 1297
rect 12371 1245 12383 1297
rect 12435 1245 12447 1297
rect 12499 1245 12511 1297
rect 12563 1282 12594 1297
rect 12563 1245 12610 1282
rect 11690 1226 12610 1245
rect 4028 1210 4294 1212
rect 6340 1041 6914 1064
rect 6340 994 6377 1041
rect 6354 989 6377 994
rect 6429 989 6441 1041
rect 6493 989 6505 1041
rect 6557 989 6569 1041
rect 6621 989 6633 1041
rect 6685 989 6697 1041
rect 6749 989 6761 1041
rect 6813 989 6825 1041
rect 6877 994 6914 1041
rect 6877 989 6900 994
rect 6354 986 6900 989
rect 3790 880 4914 964
rect 3790 658 3886 880
rect 8978 704 9034 960
rect 8960 680 9054 704
rect 3786 652 3894 658
rect 3786 618 3812 652
rect 3846 618 3894 652
rect 3786 586 3894 618
rect 8960 646 8984 680
rect 9018 646 9054 680
rect 8960 608 9054 646
rect 11674 578 12618 592
rect 11674 526 11696 578
rect 11748 526 11760 578
rect 11812 526 11824 578
rect 11876 526 11888 578
rect 11940 526 11952 578
rect 12004 526 12016 578
rect 12068 526 12080 578
rect 12132 526 12144 578
rect 12196 526 12208 578
rect 12260 526 12272 578
rect 12324 526 12336 578
rect 12388 526 12400 578
rect 12452 526 12464 578
rect 12516 526 12528 578
rect 12580 526 12618 578
rect 11674 522 12618 526
rect 3874 488 3944 494
rect 3874 436 3883 488
rect 3935 436 3944 488
rect 3874 430 3944 436
rect 9206 452 9698 472
rect 9206 400 9236 452
rect 9288 400 9300 452
rect 9352 400 9364 452
rect 9416 400 9428 452
rect 9480 400 9492 452
rect 9544 400 9556 452
rect 9608 400 9620 452
rect 9672 400 9698 452
rect 14012 428 14066 492
rect 9206 392 9698 400
<< via1 >>
rect 3872 2717 3924 2769
rect 5108 2632 5160 2684
rect 5172 2632 5224 2684
rect 5236 2632 5288 2684
rect 5300 2632 5352 2684
rect 5364 2632 5416 2684
rect 5428 2632 5480 2684
rect 5492 2632 5544 2684
rect 5556 2632 5608 2684
rect 5620 2632 5672 2684
rect 5684 2632 5736 2684
rect 5748 2632 5800 2684
rect 3874 2262 3926 2314
rect 7275 2174 7327 2226
rect 7339 2174 7391 2226
rect 7403 2174 7455 2226
rect 7467 2174 7519 2226
rect 7531 2174 7583 2226
rect 7595 2174 7647 2226
rect 7659 2174 7711 2226
rect 7723 2174 7775 2226
rect 7787 2174 7839 2226
rect 7851 2174 7903 2226
rect 5109 1878 5161 1930
rect 5173 1878 5225 1930
rect 5237 1878 5289 1930
rect 5301 1878 5353 1930
rect 5365 1878 5417 1930
rect 5429 1878 5481 1930
rect 5493 1878 5545 1930
rect 5557 1878 5609 1930
rect 5621 1878 5673 1930
rect 5685 1878 5737 1930
rect 5749 1878 5801 1930
rect 10639 1831 10691 1883
rect 10703 1831 10755 1883
rect 10767 1831 10819 1883
rect 10831 1831 10883 1883
rect 10895 1831 10947 1883
rect 10959 1831 11011 1883
rect 11023 1831 11075 1883
rect 11087 1831 11139 1883
rect 11151 1831 11203 1883
rect 11215 1831 11267 1883
rect 11279 1831 11331 1883
rect 11343 1831 11395 1883
rect 5204 1695 5256 1747
rect 5268 1695 5320 1747
rect 5332 1695 5384 1747
rect 5396 1695 5448 1747
rect 5460 1695 5512 1747
rect 5524 1695 5576 1747
rect 5588 1695 5640 1747
rect 5652 1695 5704 1747
rect 5716 1695 5768 1747
rect 5780 1695 5832 1747
rect 5844 1695 5896 1747
rect 5908 1695 5960 1747
rect 5972 1695 6024 1747
rect 6036 1695 6088 1747
rect 5168 1439 5220 1491
rect 5232 1439 5284 1491
rect 5296 1439 5348 1491
rect 5360 1439 5412 1491
rect 5424 1439 5476 1491
rect 5488 1439 5540 1491
rect 5552 1439 5604 1491
rect 5616 1439 5668 1491
rect 5680 1439 5732 1491
rect 5744 1439 5796 1491
rect 5808 1439 5860 1491
rect 5872 1439 5924 1491
rect 5936 1439 5988 1491
rect 6000 1439 6052 1491
rect 6064 1439 6116 1491
rect 6391 1384 6443 1436
rect 6455 1384 6507 1436
rect 6519 1384 6571 1436
rect 6583 1384 6635 1436
rect 6647 1384 6699 1436
rect 6711 1384 6763 1436
rect 6775 1384 6827 1436
rect 6839 1384 6891 1436
rect 10644 1432 10696 1484
rect 10708 1432 10760 1484
rect 10772 1432 10824 1484
rect 10836 1432 10888 1484
rect 10900 1432 10952 1484
rect 10964 1432 11016 1484
rect 11028 1432 11080 1484
rect 11092 1432 11144 1484
rect 11156 1432 11208 1484
rect 11220 1432 11272 1484
rect 11284 1432 11336 1484
rect 11348 1432 11400 1484
rect 7256 1304 7308 1356
rect 7320 1304 7372 1356
rect 7384 1304 7436 1356
rect 7448 1304 7500 1356
rect 7512 1304 7564 1356
rect 7576 1304 7628 1356
rect 7640 1304 7692 1356
rect 7704 1304 7756 1356
rect 7768 1304 7820 1356
rect 7832 1304 7884 1356
rect 7896 1304 7948 1356
rect 9236 1342 9288 1394
rect 9300 1342 9352 1394
rect 9364 1342 9416 1394
rect 9428 1342 9480 1394
rect 9492 1342 9544 1394
rect 9556 1342 9608 1394
rect 9620 1342 9672 1394
rect 4060 1239 4112 1291
rect 4124 1239 4176 1291
rect 4188 1239 4240 1291
rect 11743 1245 11795 1297
rect 11807 1245 11859 1297
rect 11871 1245 11923 1297
rect 11935 1245 11987 1297
rect 11999 1245 12051 1297
rect 12063 1245 12115 1297
rect 12127 1245 12179 1297
rect 12191 1245 12243 1297
rect 12255 1245 12307 1297
rect 12319 1245 12371 1297
rect 12383 1245 12435 1297
rect 12447 1245 12499 1297
rect 12511 1245 12563 1297
rect 6377 989 6429 1041
rect 6441 989 6493 1041
rect 6505 989 6557 1041
rect 6569 989 6621 1041
rect 6633 989 6685 1041
rect 6697 989 6749 1041
rect 6761 989 6813 1041
rect 6825 989 6877 1041
rect 11696 526 11748 578
rect 11760 526 11812 578
rect 11824 526 11876 578
rect 11888 526 11940 578
rect 11952 526 12004 578
rect 12016 526 12068 578
rect 12080 526 12132 578
rect 12144 526 12196 578
rect 12208 526 12260 578
rect 12272 526 12324 578
rect 12336 526 12388 578
rect 12400 526 12452 578
rect 12464 526 12516 578
rect 12528 526 12580 578
rect 3883 436 3935 488
rect 9236 400 9288 452
rect 9300 400 9352 452
rect 9364 400 9416 452
rect 9428 400 9480 452
rect 9492 400 9544 452
rect 9556 400 9608 452
rect 9620 400 9672 452
<< metal2 >>
rect 3846 2775 3940 2794
rect 3846 2719 3871 2775
rect 3927 2719 3940 2775
rect 3846 2717 3872 2719
rect 3924 2717 3940 2719
rect 3846 2686 3940 2717
rect 5092 2684 5824 2698
rect 5092 2632 5108 2684
rect 5160 2632 5172 2684
rect 5224 2632 5236 2684
rect 5288 2632 5300 2684
rect 5352 2632 5364 2684
rect 5416 2632 5428 2684
rect 5480 2632 5492 2684
rect 5544 2632 5556 2684
rect 5608 2632 5620 2684
rect 5672 2632 5684 2684
rect 5736 2632 5748 2684
rect 5800 2632 5824 2684
rect 5092 2344 5824 2632
rect 3866 2314 5824 2344
rect 3866 2262 3874 2314
rect 3926 2262 5824 2314
rect 3866 2226 5824 2262
rect 3954 2220 5824 2226
rect 5092 1930 5824 2220
rect 5092 1878 5109 1930
rect 5161 1878 5173 1930
rect 5225 1878 5237 1930
rect 5289 1878 5301 1930
rect 5353 1878 5365 1930
rect 5417 1878 5429 1930
rect 5481 1878 5493 1930
rect 5545 1878 5557 1930
rect 5609 1878 5621 1930
rect 5673 1878 5685 1930
rect 5737 1878 5749 1930
rect 5801 1878 5824 1930
rect 5092 1870 5824 1878
rect 7214 2226 7992 2234
rect 7214 2174 7275 2226
rect 7327 2174 7339 2226
rect 7391 2174 7403 2226
rect 7455 2174 7467 2226
rect 7519 2174 7531 2226
rect 7583 2174 7595 2226
rect 7647 2174 7659 2226
rect 7711 2174 7723 2226
rect 7775 2174 7787 2226
rect 7839 2174 7851 2226
rect 7903 2174 7992 2226
rect 5160 1747 6130 1772
rect 5160 1695 5204 1747
rect 5256 1695 5268 1747
rect 5320 1695 5332 1747
rect 5384 1695 5396 1747
rect 5448 1695 5460 1747
rect 5512 1695 5524 1747
rect 5576 1695 5588 1747
rect 5640 1695 5652 1747
rect 5704 1695 5716 1747
rect 5768 1695 5780 1747
rect 5832 1695 5844 1747
rect 5896 1695 5908 1747
rect 5960 1695 5972 1747
rect 6024 1695 6036 1747
rect 6088 1695 6130 1747
rect 5160 1542 6130 1695
rect 5164 1491 6130 1542
rect 5164 1439 5168 1491
rect 5220 1439 5232 1491
rect 5284 1439 5296 1491
rect 5348 1439 5360 1491
rect 5412 1439 5424 1491
rect 5476 1439 5488 1491
rect 5540 1439 5552 1491
rect 5604 1439 5616 1491
rect 5668 1439 5680 1491
rect 5732 1439 5744 1491
rect 5796 1439 5808 1491
rect 5860 1439 5872 1491
rect 5924 1439 5936 1491
rect 5988 1439 6000 1491
rect 6052 1439 6064 1491
rect 6116 1439 6130 1491
rect 5164 1418 6130 1439
rect 6338 1436 6932 1444
rect 5164 1394 5326 1418
rect 6338 1384 6391 1436
rect 6443 1384 6455 1436
rect 6507 1384 6519 1436
rect 6571 1384 6583 1436
rect 6635 1384 6647 1436
rect 6699 1384 6711 1436
rect 6763 1384 6775 1436
rect 6827 1384 6839 1436
rect 6891 1384 6932 1436
rect 3954 1326 4292 1330
rect 3866 1299 4292 1326
rect 3866 1243 3886 1299
rect 3942 1291 4292 1299
rect 3942 1243 4060 1291
rect 3866 1239 4060 1243
rect 4112 1239 4124 1291
rect 4176 1239 4188 1291
rect 4240 1239 4292 1291
rect 3866 1210 4292 1239
rect 3870 494 3936 1210
rect 6338 1041 6932 1384
rect 7214 1356 7992 2174
rect 10606 1883 11466 1896
rect 10606 1831 10639 1883
rect 10691 1831 10703 1883
rect 10755 1831 10767 1883
rect 10819 1831 10831 1883
rect 10883 1831 10895 1883
rect 10947 1831 10959 1883
rect 11011 1831 11023 1883
rect 11075 1831 11087 1883
rect 11139 1831 11151 1883
rect 11203 1831 11215 1883
rect 11267 1831 11279 1883
rect 11331 1831 11343 1883
rect 11395 1831 11466 1883
rect 10606 1484 11466 1831
rect 10606 1432 10644 1484
rect 10696 1432 10708 1484
rect 10760 1432 10772 1484
rect 10824 1432 10836 1484
rect 10888 1432 10900 1484
rect 10952 1432 10964 1484
rect 11016 1432 11028 1484
rect 11080 1432 11092 1484
rect 11144 1432 11156 1484
rect 11208 1432 11220 1484
rect 11272 1432 11284 1484
rect 11336 1432 11348 1484
rect 11400 1432 11466 1484
rect 10606 1420 11466 1432
rect 7214 1304 7256 1356
rect 7308 1304 7320 1356
rect 7372 1304 7384 1356
rect 7436 1304 7448 1356
rect 7500 1304 7512 1356
rect 7564 1304 7576 1356
rect 7628 1304 7640 1356
rect 7692 1304 7704 1356
rect 7756 1304 7768 1356
rect 7820 1304 7832 1356
rect 7884 1304 7896 1356
rect 7948 1304 7992 1356
rect 7214 1290 7992 1304
rect 9206 1394 9706 1404
rect 9206 1342 9236 1394
rect 9288 1342 9300 1394
rect 9352 1342 9364 1394
rect 9416 1342 9428 1394
rect 9480 1342 9492 1394
rect 9544 1342 9556 1394
rect 9608 1342 9620 1394
rect 9672 1342 9706 1394
rect 6338 989 6377 1041
rect 6429 989 6441 1041
rect 6493 989 6505 1041
rect 6557 989 6569 1041
rect 6621 989 6633 1041
rect 6685 989 6697 1041
rect 6749 989 6761 1041
rect 6813 989 6825 1041
rect 6877 989 6932 1041
rect 6338 980 6932 989
rect 9206 598 9706 1342
rect 3870 488 3944 494
rect 3870 436 3883 488
rect 3935 436 3944 488
rect 3870 430 3944 436
rect 9204 452 9706 598
rect 11684 1297 12628 1312
rect 11684 1245 11743 1297
rect 11795 1245 11807 1297
rect 11859 1245 11871 1297
rect 11923 1245 11935 1297
rect 11987 1245 11999 1297
rect 12051 1245 12063 1297
rect 12115 1245 12127 1297
rect 12179 1245 12191 1297
rect 12243 1245 12255 1297
rect 12307 1245 12319 1297
rect 12371 1245 12383 1297
rect 12435 1245 12447 1297
rect 12499 1245 12511 1297
rect 12563 1245 12628 1297
rect 11684 578 12628 1245
rect 11684 526 11696 578
rect 11748 526 11760 578
rect 11812 526 11824 578
rect 11876 526 11888 578
rect 11940 526 11952 578
rect 12004 526 12016 578
rect 12068 526 12080 578
rect 12132 526 12144 578
rect 12196 526 12208 578
rect 12260 526 12272 578
rect 12324 526 12336 578
rect 12388 526 12400 578
rect 12452 526 12464 578
rect 12516 526 12528 578
rect 12580 526 12628 578
rect 11684 514 12628 526
rect 9204 400 9236 452
rect 9288 400 9300 452
rect 9352 400 9364 452
rect 9416 400 9428 452
rect 9480 400 9492 452
rect 9544 400 9556 452
rect 9608 400 9620 452
rect 9672 400 9706 452
rect 9204 386 9706 400
rect 9204 -276 9704 386
<< via2 >>
rect 3871 2769 3927 2775
rect 3871 2719 3872 2769
rect 3872 2719 3924 2769
rect 3924 2719 3927 2769
rect 3886 1243 3942 1299
<< metal3 >>
rect 3836 2775 3950 2804
rect 3836 2719 3871 2775
rect 3927 2719 3950 2775
rect 3836 2668 3950 2719
rect 3878 1299 3948 2668
rect 3878 1243 3886 1299
rect 3942 1243 3948 1299
rect 3878 1208 3948 1243
use sky130_fd_pr__nfet_01v8_lvt_8K7EBA  sky130_fd_pr__nfet_01v8_lvt_8K7EBA_0
timestamp 1640969486
transform 0 1 6946 -1 0 925
box -221 -2200 221 2200
use sky130_fd_pr__nfet_01v8_lvt_8K7EBA  sky130_fd_pr__nfet_01v8_lvt_8K7EBA_1
timestamp 1640969486
transform 0 -1 6946 -1 0 1369
box -221 -2200 221 2200
use sky130_fd_pr__nfet_01v8_lvt_8K7EBA  sky130_fd_pr__nfet_01v8_lvt_8K7EBA_2
timestamp 1640969486
transform 0 1 6946 -1 0 1823
box -221 -2200 221 2200
use sky130_fd_pr__nfet_01v8_lvt_8K7EBA  sky130_fd_pr__nfet_01v8_lvt_8K7EBA_3
timestamp 1640969486
transform 0 1 11980 -1 0 1367
box -221 -2200 221 2200
use sky130_fd_pr__nfet_01v8_lvt_8K7EBA  sky130_fd_pr__nfet_01v8_lvt_8K7EBA_4
timestamp 1640969486
transform 0 1 11980 -1 0 1825
box -221 -2200 221 2200
use sky130_fd_pr__pfet_01v8_lvt_4QC8GG  sky130_fd_pr__pfet_01v8_lvt_4QC8GG_0
timestamp 1640969486
transform 0 1 8971 -1 0 2287
box -231 -5219 231 5219
use sky130_fd_pr__pfet_01v8_lvt_4QC8GG  sky130_fd_pr__pfet_01v8_lvt_4QC8GG_1
timestamp 1640969486
transform 0 1 8971 -1 0 2745
box -231 -5219 231 5219
use sky130_fd_pr__pfet_01v8_lvt_4QC8GG  sky130_fd_pr__pfet_01v8_lvt_4QC8GG_2
timestamp 1640969486
transform 0 1 8973 -1 0 459
box -231 -5219 231 5219
<< labels >>
rlabel metal1 s 3816 1492 3816 1492 4 VIN-
port 1 nsew
rlabel metal2 s 12062 882 12062 882 4 VOUT
port 2 nsew
rlabel locali s 14138 1550 14138 1550 4 VSS
port 3 nsew
rlabel metal2 s 9454 -218 9454 -218 4 VINp
port 4 nsew
<< end >>
