magic
tech sky130A
magscale 1 2
timestamp 1640969486
<< pwell >>
rect -134 -1076 134 1076
<< nmos >>
rect -50 -1050 50 1050
<< ndiff >>
rect -108 1037 -50 1050
rect -108 1003 -96 1037
rect -62 1003 -50 1037
rect -108 969 -50 1003
rect -108 935 -96 969
rect -62 935 -50 969
rect -108 901 -50 935
rect -108 867 -96 901
rect -62 867 -50 901
rect -108 833 -50 867
rect -108 799 -96 833
rect -62 799 -50 833
rect -108 765 -50 799
rect -108 731 -96 765
rect -62 731 -50 765
rect -108 697 -50 731
rect -108 663 -96 697
rect -62 663 -50 697
rect -108 629 -50 663
rect -108 595 -96 629
rect -62 595 -50 629
rect -108 561 -50 595
rect -108 527 -96 561
rect -62 527 -50 561
rect -108 493 -50 527
rect -108 459 -96 493
rect -62 459 -50 493
rect -108 425 -50 459
rect -108 391 -96 425
rect -62 391 -50 425
rect -108 357 -50 391
rect -108 323 -96 357
rect -62 323 -50 357
rect -108 289 -50 323
rect -108 255 -96 289
rect -62 255 -50 289
rect -108 221 -50 255
rect -108 187 -96 221
rect -62 187 -50 221
rect -108 153 -50 187
rect -108 119 -96 153
rect -62 119 -50 153
rect -108 85 -50 119
rect -108 51 -96 85
rect -62 51 -50 85
rect -108 17 -50 51
rect -108 -17 -96 17
rect -62 -17 -50 17
rect -108 -51 -50 -17
rect -108 -85 -96 -51
rect -62 -85 -50 -51
rect -108 -119 -50 -85
rect -108 -153 -96 -119
rect -62 -153 -50 -119
rect -108 -187 -50 -153
rect -108 -221 -96 -187
rect -62 -221 -50 -187
rect -108 -255 -50 -221
rect -108 -289 -96 -255
rect -62 -289 -50 -255
rect -108 -323 -50 -289
rect -108 -357 -96 -323
rect -62 -357 -50 -323
rect -108 -391 -50 -357
rect -108 -425 -96 -391
rect -62 -425 -50 -391
rect -108 -459 -50 -425
rect -108 -493 -96 -459
rect -62 -493 -50 -459
rect -108 -527 -50 -493
rect -108 -561 -96 -527
rect -62 -561 -50 -527
rect -108 -595 -50 -561
rect -108 -629 -96 -595
rect -62 -629 -50 -595
rect -108 -663 -50 -629
rect -108 -697 -96 -663
rect -62 -697 -50 -663
rect -108 -731 -50 -697
rect -108 -765 -96 -731
rect -62 -765 -50 -731
rect -108 -799 -50 -765
rect -108 -833 -96 -799
rect -62 -833 -50 -799
rect -108 -867 -50 -833
rect -108 -901 -96 -867
rect -62 -901 -50 -867
rect -108 -935 -50 -901
rect -108 -969 -96 -935
rect -62 -969 -50 -935
rect -108 -1003 -50 -969
rect -108 -1037 -96 -1003
rect -62 -1037 -50 -1003
rect -108 -1050 -50 -1037
rect 50 1037 108 1050
rect 50 1003 62 1037
rect 96 1003 108 1037
rect 50 969 108 1003
rect 50 935 62 969
rect 96 935 108 969
rect 50 901 108 935
rect 50 867 62 901
rect 96 867 108 901
rect 50 833 108 867
rect 50 799 62 833
rect 96 799 108 833
rect 50 765 108 799
rect 50 731 62 765
rect 96 731 108 765
rect 50 697 108 731
rect 50 663 62 697
rect 96 663 108 697
rect 50 629 108 663
rect 50 595 62 629
rect 96 595 108 629
rect 50 561 108 595
rect 50 527 62 561
rect 96 527 108 561
rect 50 493 108 527
rect 50 459 62 493
rect 96 459 108 493
rect 50 425 108 459
rect 50 391 62 425
rect 96 391 108 425
rect 50 357 108 391
rect 50 323 62 357
rect 96 323 108 357
rect 50 289 108 323
rect 50 255 62 289
rect 96 255 108 289
rect 50 221 108 255
rect 50 187 62 221
rect 96 187 108 221
rect 50 153 108 187
rect 50 119 62 153
rect 96 119 108 153
rect 50 85 108 119
rect 50 51 62 85
rect 96 51 108 85
rect 50 17 108 51
rect 50 -17 62 17
rect 96 -17 108 17
rect 50 -51 108 -17
rect 50 -85 62 -51
rect 96 -85 108 -51
rect 50 -119 108 -85
rect 50 -153 62 -119
rect 96 -153 108 -119
rect 50 -187 108 -153
rect 50 -221 62 -187
rect 96 -221 108 -187
rect 50 -255 108 -221
rect 50 -289 62 -255
rect 96 -289 108 -255
rect 50 -323 108 -289
rect 50 -357 62 -323
rect 96 -357 108 -323
rect 50 -391 108 -357
rect 50 -425 62 -391
rect 96 -425 108 -391
rect 50 -459 108 -425
rect 50 -493 62 -459
rect 96 -493 108 -459
rect 50 -527 108 -493
rect 50 -561 62 -527
rect 96 -561 108 -527
rect 50 -595 108 -561
rect 50 -629 62 -595
rect 96 -629 108 -595
rect 50 -663 108 -629
rect 50 -697 62 -663
rect 96 -697 108 -663
rect 50 -731 108 -697
rect 50 -765 62 -731
rect 96 -765 108 -731
rect 50 -799 108 -765
rect 50 -833 62 -799
rect 96 -833 108 -799
rect 50 -867 108 -833
rect 50 -901 62 -867
rect 96 -901 108 -867
rect 50 -935 108 -901
rect 50 -969 62 -935
rect 96 -969 108 -935
rect 50 -1003 108 -969
rect 50 -1037 62 -1003
rect 96 -1037 108 -1003
rect 50 -1050 108 -1037
<< ndiffc >>
rect -96 1003 -62 1037
rect -96 935 -62 969
rect -96 867 -62 901
rect -96 799 -62 833
rect -96 731 -62 765
rect -96 663 -62 697
rect -96 595 -62 629
rect -96 527 -62 561
rect -96 459 -62 493
rect -96 391 -62 425
rect -96 323 -62 357
rect -96 255 -62 289
rect -96 187 -62 221
rect -96 119 -62 153
rect -96 51 -62 85
rect -96 -17 -62 17
rect -96 -85 -62 -51
rect -96 -153 -62 -119
rect -96 -221 -62 -187
rect -96 -289 -62 -255
rect -96 -357 -62 -323
rect -96 -425 -62 -391
rect -96 -493 -62 -459
rect -96 -561 -62 -527
rect -96 -629 -62 -595
rect -96 -697 -62 -663
rect -96 -765 -62 -731
rect -96 -833 -62 -799
rect -96 -901 -62 -867
rect -96 -969 -62 -935
rect -96 -1037 -62 -1003
rect 62 1003 96 1037
rect 62 935 96 969
rect 62 867 96 901
rect 62 799 96 833
rect 62 731 96 765
rect 62 663 96 697
rect 62 595 96 629
rect 62 527 96 561
rect 62 459 96 493
rect 62 391 96 425
rect 62 323 96 357
rect 62 255 96 289
rect 62 187 96 221
rect 62 119 96 153
rect 62 51 96 85
rect 62 -17 96 17
rect 62 -85 96 -51
rect 62 -153 96 -119
rect 62 -221 96 -187
rect 62 -289 96 -255
rect 62 -357 96 -323
rect 62 -425 96 -391
rect 62 -493 96 -459
rect 62 -561 96 -527
rect 62 -629 96 -595
rect 62 -697 96 -663
rect 62 -765 96 -731
rect 62 -833 96 -799
rect 62 -901 96 -867
rect 62 -969 96 -935
rect 62 -1037 96 -1003
<< poly >>
rect -50 1050 50 1076
rect -50 -1076 50 -1050
<< locali >>
rect -96 1037 -62 1054
rect -96 969 -62 991
rect -96 901 -62 919
rect -96 833 -62 847
rect -96 765 -62 775
rect -96 697 -62 703
rect -96 629 -62 631
rect -96 593 -62 595
rect -96 521 -62 527
rect -96 449 -62 459
rect -96 377 -62 391
rect -96 305 -62 323
rect -96 233 -62 255
rect -96 161 -62 187
rect -96 89 -62 119
rect -96 17 -62 51
rect -96 -51 -62 -17
rect -96 -119 -62 -89
rect -96 -187 -62 -161
rect -96 -255 -62 -233
rect -96 -323 -62 -305
rect -96 -391 -62 -377
rect -96 -459 -62 -449
rect -96 -527 -62 -521
rect -96 -595 -62 -593
rect -96 -631 -62 -629
rect -96 -703 -62 -697
rect -96 -775 -62 -765
rect -96 -847 -62 -833
rect -96 -919 -62 -901
rect -96 -991 -62 -969
rect -96 -1054 -62 -1037
rect 62 1037 96 1054
rect 62 969 96 991
rect 62 901 96 919
rect 62 833 96 847
rect 62 765 96 775
rect 62 697 96 703
rect 62 629 96 631
rect 62 593 96 595
rect 62 521 96 527
rect 62 449 96 459
rect 62 377 96 391
rect 62 305 96 323
rect 62 233 96 255
rect 62 161 96 187
rect 62 89 96 119
rect 62 17 96 51
rect 62 -51 96 -17
rect 62 -119 96 -89
rect 62 -187 96 -161
rect 62 -255 96 -233
rect 62 -323 96 -305
rect 62 -391 96 -377
rect 62 -459 96 -449
rect 62 -527 96 -521
rect 62 -595 96 -593
rect 62 -631 96 -629
rect 62 -703 96 -697
rect 62 -775 96 -765
rect 62 -847 96 -833
rect 62 -919 96 -901
rect 62 -991 96 -969
rect 62 -1054 96 -1037
<< viali >>
rect -96 1003 -62 1025
rect -96 991 -62 1003
rect -96 935 -62 953
rect -96 919 -62 935
rect -96 867 -62 881
rect -96 847 -62 867
rect -96 799 -62 809
rect -96 775 -62 799
rect -96 731 -62 737
rect -96 703 -62 731
rect -96 663 -62 665
rect -96 631 -62 663
rect -96 561 -62 593
rect -96 559 -62 561
rect -96 493 -62 521
rect -96 487 -62 493
rect -96 425 -62 449
rect -96 415 -62 425
rect -96 357 -62 377
rect -96 343 -62 357
rect -96 289 -62 305
rect -96 271 -62 289
rect -96 221 -62 233
rect -96 199 -62 221
rect -96 153 -62 161
rect -96 127 -62 153
rect -96 85 -62 89
rect -96 55 -62 85
rect -96 -17 -62 17
rect -96 -85 -62 -55
rect -96 -89 -62 -85
rect -96 -153 -62 -127
rect -96 -161 -62 -153
rect -96 -221 -62 -199
rect -96 -233 -62 -221
rect -96 -289 -62 -271
rect -96 -305 -62 -289
rect -96 -357 -62 -343
rect -96 -377 -62 -357
rect -96 -425 -62 -415
rect -96 -449 -62 -425
rect -96 -493 -62 -487
rect -96 -521 -62 -493
rect -96 -561 -62 -559
rect -96 -593 -62 -561
rect -96 -663 -62 -631
rect -96 -665 -62 -663
rect -96 -731 -62 -703
rect -96 -737 -62 -731
rect -96 -799 -62 -775
rect -96 -809 -62 -799
rect -96 -867 -62 -847
rect -96 -881 -62 -867
rect -96 -935 -62 -919
rect -96 -953 -62 -935
rect -96 -1003 -62 -991
rect -96 -1025 -62 -1003
rect 62 1003 96 1025
rect 62 991 96 1003
rect 62 935 96 953
rect 62 919 96 935
rect 62 867 96 881
rect 62 847 96 867
rect 62 799 96 809
rect 62 775 96 799
rect 62 731 96 737
rect 62 703 96 731
rect 62 663 96 665
rect 62 631 96 663
rect 62 561 96 593
rect 62 559 96 561
rect 62 493 96 521
rect 62 487 96 493
rect 62 425 96 449
rect 62 415 96 425
rect 62 357 96 377
rect 62 343 96 357
rect 62 289 96 305
rect 62 271 96 289
rect 62 221 96 233
rect 62 199 96 221
rect 62 153 96 161
rect 62 127 96 153
rect 62 85 96 89
rect 62 55 96 85
rect 62 -17 96 17
rect 62 -85 96 -55
rect 62 -89 96 -85
rect 62 -153 96 -127
rect 62 -161 96 -153
rect 62 -221 96 -199
rect 62 -233 96 -221
rect 62 -289 96 -271
rect 62 -305 96 -289
rect 62 -357 96 -343
rect 62 -377 96 -357
rect 62 -425 96 -415
rect 62 -449 96 -425
rect 62 -493 96 -487
rect 62 -521 96 -493
rect 62 -561 96 -559
rect 62 -593 96 -561
rect 62 -663 96 -631
rect 62 -665 96 -663
rect 62 -731 96 -703
rect 62 -737 96 -731
rect 62 -799 96 -775
rect 62 -809 96 -799
rect 62 -867 96 -847
rect 62 -881 96 -867
rect 62 -935 96 -919
rect 62 -953 96 -935
rect 62 -1003 96 -991
rect 62 -1025 96 -1003
<< metal1 >>
rect -102 1025 -56 1050
rect -102 991 -96 1025
rect -62 991 -56 1025
rect -102 953 -56 991
rect -102 919 -96 953
rect -62 919 -56 953
rect -102 881 -56 919
rect -102 847 -96 881
rect -62 847 -56 881
rect -102 809 -56 847
rect -102 775 -96 809
rect -62 775 -56 809
rect -102 737 -56 775
rect -102 703 -96 737
rect -62 703 -56 737
rect -102 665 -56 703
rect -102 631 -96 665
rect -62 631 -56 665
rect -102 593 -56 631
rect -102 559 -96 593
rect -62 559 -56 593
rect -102 521 -56 559
rect -102 487 -96 521
rect -62 487 -56 521
rect -102 449 -56 487
rect -102 415 -96 449
rect -62 415 -56 449
rect -102 377 -56 415
rect -102 343 -96 377
rect -62 343 -56 377
rect -102 305 -56 343
rect -102 271 -96 305
rect -62 271 -56 305
rect -102 233 -56 271
rect -102 199 -96 233
rect -62 199 -56 233
rect -102 161 -56 199
rect -102 127 -96 161
rect -62 127 -56 161
rect -102 89 -56 127
rect -102 55 -96 89
rect -62 55 -56 89
rect -102 17 -56 55
rect -102 -17 -96 17
rect -62 -17 -56 17
rect -102 -55 -56 -17
rect -102 -89 -96 -55
rect -62 -89 -56 -55
rect -102 -127 -56 -89
rect -102 -161 -96 -127
rect -62 -161 -56 -127
rect -102 -199 -56 -161
rect -102 -233 -96 -199
rect -62 -233 -56 -199
rect -102 -271 -56 -233
rect -102 -305 -96 -271
rect -62 -305 -56 -271
rect -102 -343 -56 -305
rect -102 -377 -96 -343
rect -62 -377 -56 -343
rect -102 -415 -56 -377
rect -102 -449 -96 -415
rect -62 -449 -56 -415
rect -102 -487 -56 -449
rect -102 -521 -96 -487
rect -62 -521 -56 -487
rect -102 -559 -56 -521
rect -102 -593 -96 -559
rect -62 -593 -56 -559
rect -102 -631 -56 -593
rect -102 -665 -96 -631
rect -62 -665 -56 -631
rect -102 -703 -56 -665
rect -102 -737 -96 -703
rect -62 -737 -56 -703
rect -102 -775 -56 -737
rect -102 -809 -96 -775
rect -62 -809 -56 -775
rect -102 -847 -56 -809
rect -102 -881 -96 -847
rect -62 -881 -56 -847
rect -102 -919 -56 -881
rect -102 -953 -96 -919
rect -62 -953 -56 -919
rect -102 -991 -56 -953
rect -102 -1025 -96 -991
rect -62 -1025 -56 -991
rect -102 -1050 -56 -1025
rect 56 1025 102 1050
rect 56 991 62 1025
rect 96 991 102 1025
rect 56 953 102 991
rect 56 919 62 953
rect 96 919 102 953
rect 56 881 102 919
rect 56 847 62 881
rect 96 847 102 881
rect 56 809 102 847
rect 56 775 62 809
rect 96 775 102 809
rect 56 737 102 775
rect 56 703 62 737
rect 96 703 102 737
rect 56 665 102 703
rect 56 631 62 665
rect 96 631 102 665
rect 56 593 102 631
rect 56 559 62 593
rect 96 559 102 593
rect 56 521 102 559
rect 56 487 62 521
rect 96 487 102 521
rect 56 449 102 487
rect 56 415 62 449
rect 96 415 102 449
rect 56 377 102 415
rect 56 343 62 377
rect 96 343 102 377
rect 56 305 102 343
rect 56 271 62 305
rect 96 271 102 305
rect 56 233 102 271
rect 56 199 62 233
rect 96 199 102 233
rect 56 161 102 199
rect 56 127 62 161
rect 96 127 102 161
rect 56 89 102 127
rect 56 55 62 89
rect 96 55 102 89
rect 56 17 102 55
rect 56 -17 62 17
rect 96 -17 102 17
rect 56 -55 102 -17
rect 56 -89 62 -55
rect 96 -89 102 -55
rect 56 -127 102 -89
rect 56 -161 62 -127
rect 96 -161 102 -127
rect 56 -199 102 -161
rect 56 -233 62 -199
rect 96 -233 102 -199
rect 56 -271 102 -233
rect 56 -305 62 -271
rect 96 -305 102 -271
rect 56 -343 102 -305
rect 56 -377 62 -343
rect 96 -377 102 -343
rect 56 -415 102 -377
rect 56 -449 62 -415
rect 96 -449 102 -415
rect 56 -487 102 -449
rect 56 -521 62 -487
rect 96 -521 102 -487
rect 56 -559 102 -521
rect 56 -593 62 -559
rect 96 -593 102 -559
rect 56 -631 102 -593
rect 56 -665 62 -631
rect 96 -665 102 -631
rect 56 -703 102 -665
rect 56 -737 62 -703
rect 96 -737 102 -703
rect 56 -775 102 -737
rect 56 -809 62 -775
rect 96 -809 102 -775
rect 56 -847 102 -809
rect 56 -881 62 -847
rect 96 -881 102 -847
rect 56 -919 102 -881
rect 56 -953 62 -919
rect 96 -953 102 -919
rect 56 -991 102 -953
rect 56 -1025 62 -991
rect 96 -1025 102 -991
rect 56 -1050 102 -1025
<< end >>
