magic
tech sky130A
magscale 1 2
timestamp 1640969486
<< metal1 >>
rect -480 38310 948 38438
rect -480 37938 -281 38310
rect 539 37938 948 38310
rect -480 37872 948 37938
rect -480 37868 -396 37872
rect 848 37792 948 37872
rect 882 37746 948 37792
rect 882 37730 904 37746
rect 936 37556 948 37746
rect 17684 520 18170 594
rect 17684 514 18210 520
rect 17435 423 18210 514
rect 17435 179 17843 423
rect 18087 179 18210 423
rect 17435 56 18210 179
rect 17714 42 18210 56
<< via1 >>
rect -281 37938 539 38310
rect 17843 179 18087 423
<< metal2 >>
rect -390 39892 590 40110
rect -390 39196 -256 39892
rect 440 39196 590 39892
rect -390 38592 590 39196
rect -396 38310 660 38592
rect -396 37938 -281 38310
rect 539 37938 660 38310
rect -396 37894 660 37938
rect -390 37890 -246 37894
rect 480 37890 590 37894
rect 17714 423 18210 520
rect 17714 179 17843 423
rect 18087 179 18210 423
rect 17714 42 18210 179
rect 17770 30 18164 42
<< via2 >>
rect -256 39196 440 39892
rect 17857 193 18073 409
<< metal3 >>
rect -390 39892 624 45240
rect -390 39196 -256 39892
rect 440 39196 624 39892
rect -390 38960 624 39196
rect 17714 413 18210 520
rect 17714 189 17853 413
rect 18077 189 18210 413
rect 17714 42 18210 189
rect 17770 30 18164 42
<< via3 >>
rect 17853 409 18077 413
rect 17853 193 17857 409
rect 17857 193 18073 409
rect 18073 193 18077 409
rect 17853 189 18077 193
<< metal4 >>
rect 14870 40532 16038 44810
rect 14870 40064 18172 40532
rect 17760 520 18152 40064
rect 17714 413 18210 520
rect 17714 189 17853 413
rect 18077 189 18210 413
rect 17714 42 18210 189
use FINAL  FINAL_0
timestamp 1640969486
transform 1 0 2 0 1 2
box -2 -2 136810 98784
use cap_30_layout  cap_30_layout_0
timestamp 1640969486
transform 1 0 12438 0 1 62996
box -19594 -20254 7036 8558
<< labels >>
rlabel metal3 s 326 40778 326 40778 4 VINN
port 1 nsew
rlabel metal2 s -72 38660 -72 38660 4 VINN
port 1 nsew
rlabel metal4 s 17974 40444 17974 40444 4 VINP
port 2 nsew
<< end >>
