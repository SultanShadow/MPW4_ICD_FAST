magic
tech sky130A
magscale 1 2
timestamp 1640969486
<< nwell >>
rect 4753 3005 4825 3075
rect 4929 3005 5001 3075
rect 5105 3005 5177 3075
rect 5281 3005 5353 3075
rect 5457 3005 5529 3075
<< locali >>
rect 4577 3057 4649 3075
rect 4577 3023 4596 3057
rect 4630 3023 4649 3057
rect 4577 3005 4649 3023
rect 4753 3057 4825 3075
rect 4753 3023 4772 3057
rect 4806 3023 4825 3057
rect 4753 3005 4825 3023
rect 4929 3057 5001 3075
rect 4929 3023 4948 3057
rect 4982 3023 5001 3057
rect 4929 3005 5001 3023
rect 5105 3057 5177 3075
rect 5105 3023 5124 3057
rect 5158 3023 5177 3057
rect 5105 3005 5177 3023
rect 5281 3057 5353 3075
rect 5281 3023 5300 3057
rect 5334 3023 5353 3057
rect 5281 3005 5353 3023
rect 5457 3057 5529 3075
rect 5457 3023 5476 3057
rect 5510 3023 5529 3057
rect 5457 3005 5529 3023
rect 834 -382 2630 283
rect 8 -840 2630 -382
rect 834 -1005 2630 -840
rect 2980 -995 3930 310
rect 566 -1304 736 -1028
rect 959 -1299 1759 -1287
rect 86 -1553 101 -1519
rect 135 -1553 173 -1519
rect 207 -1553 245 -1519
rect 279 -1553 295 -1519
rect 959 -1630 1990 -1299
rect 2961 -1319 4376 -1174
rect 959 -1648 1759 -1630
rect 849 -1927 1640 -1910
rect 474 -2476 594 -2144
rect 849 -2169 1986 -1927
rect 849 -2179 1640 -2169
<< viali >>
rect 4596 3023 4630 3057
rect 4772 3023 4806 3057
rect 4948 3023 4982 3057
rect 5124 3023 5158 3057
rect 5300 3023 5334 3057
rect 5476 3023 5510 3057
rect 101 -1553 135 -1519
rect 173 -1553 207 -1519
rect 245 -1553 279 -1519
<< metal1 >>
rect 5598 5234 6094 5235
rect 1501 5213 6094 5234
rect 1501 5212 5630 5213
rect 1501 4904 4591 5212
rect 5475 4905 5630 5212
rect 6066 4905 6094 5213
rect 5475 4904 6094 4905
rect 1501 4885 6094 4904
rect 535 3968 1497 4011
rect 535 3724 571 3968
rect 1007 3724 1497 3968
rect 535 3674 1497 3724
rect 4577 3065 5529 3075
rect 4577 3013 4587 3065
rect 4639 3013 4763 3065
rect 4815 3013 4939 3065
rect 4991 3013 5115 3065
rect 5167 3013 5291 3065
rect 5343 3013 5467 3065
rect 5519 3013 5529 3065
rect 2228 3008 2232 3010
rect 4577 3005 5529 3013
rect 5603 2711 6094 2721
rect 5603 2659 5630 2711
rect 5682 2659 5694 2711
rect 5746 2659 5758 2711
rect 5810 2659 5822 2711
rect 5874 2659 5886 2711
rect 5938 2659 5950 2711
rect 6002 2659 6014 2711
rect 6066 2659 6094 2711
rect 5603 2651 6094 2659
rect 0 583 17 705
rect -646 -603 -96 -486
rect -646 -2511 -452 -603
rect -208 -1113 -96 -603
rect 1279 -1012 1727 498
rect 2064 -1012 2512 503
rect 2968 -1012 3416 535
rect 3709 -1012 4157 507
rect 880 -1073 4407 -1012
rect -208 -1179 848 -1113
rect 880 -1119 2480 -1073
rect -208 -2275 -96 -1179
rect 56 -1519 314 -1490
rect 56 -1553 101 -1519
rect 135 -1553 173 -1519
rect 207 -1553 245 -1519
rect 279 -1553 314 -1519
rect 56 -1970 314 -1553
rect 949 -1814 1381 -1178
rect 2512 -1179 2568 -1113
rect 2864 -1179 2920 -1113
rect 2952 -1119 4407 -1073
rect 4464 -1179 4671 -1113
rect 2161 -1744 2442 -1742
rect 1480 -1754 6094 -1744
rect 1480 -1806 5631 -1754
rect 5683 -1806 5695 -1754
rect 5747 -1806 5759 -1754
rect 5811 -1806 5823 -1754
rect 5875 -1806 5887 -1754
rect 5939 -1806 5951 -1754
rect 6003 -1806 6015 -1754
rect 6067 -1806 6094 -1754
rect 1480 -1814 6094 -1806
rect 2161 -1970 2442 -1814
rect 56 -2196 2442 -1970
rect -208 -2345 1134 -2275
rect 3134 -2345 3743 -2275
rect -208 -2511 -96 -2345
rect -646 -2615 -96 -2511
<< via1 >>
rect 4591 4904 5475 5212
rect 5630 4905 6066 5213
rect 571 3724 1007 3968
rect 4587 3057 4639 3065
rect 4587 3023 4596 3057
rect 4596 3023 4630 3057
rect 4630 3023 4639 3057
rect 4587 3013 4639 3023
rect 4763 3057 4815 3065
rect 4763 3023 4772 3057
rect 4772 3023 4806 3057
rect 4806 3023 4815 3057
rect 4763 3013 4815 3023
rect 4939 3057 4991 3065
rect 4939 3023 4948 3057
rect 4948 3023 4982 3057
rect 4982 3023 4991 3057
rect 4939 3013 4991 3023
rect 5115 3057 5167 3065
rect 5115 3023 5124 3057
rect 5124 3023 5158 3057
rect 5158 3023 5167 3057
rect 5115 3013 5167 3023
rect 5291 3057 5343 3065
rect 5291 3023 5300 3057
rect 5300 3023 5334 3057
rect 5334 3023 5343 3057
rect 5291 3013 5343 3023
rect 5467 3057 5519 3065
rect 5467 3023 5476 3057
rect 5476 3023 5510 3057
rect 5510 3023 5519 3057
rect 5467 3013 5519 3023
rect 5630 2659 5682 2711
rect 5694 2659 5746 2711
rect 5758 2659 5810 2711
rect 5822 2659 5874 2711
rect 5886 2659 5938 2711
rect 5950 2659 6002 2711
rect 6014 2659 6066 2711
rect -452 -2511 -208 -603
rect 5631 -1806 5683 -1754
rect 5695 -1806 5747 -1754
rect 5759 -1806 5811 -1754
rect 5823 -1806 5875 -1754
rect 5887 -1806 5939 -1754
rect 5951 -1806 6003 -1754
rect 6015 -1806 6067 -1754
<< metal2 >>
rect 4577 5213 6094 5235
rect 4577 5212 5630 5213
rect 4577 4904 4591 5212
rect 5475 4905 5630 5212
rect 6066 4905 6094 5213
rect 5475 4904 6094 4905
rect -90 3968 1069 4006
rect -90 3947 571 3968
rect -90 3731 -49 3947
rect 407 3731 571 3947
rect -90 3724 571 3731
rect 1007 3724 1069 3968
rect -90 3674 1069 3724
rect 4577 3065 6094 4904
rect 4577 3013 4587 3065
rect 4639 3013 4763 3065
rect 4815 3013 4939 3065
rect 4991 3013 5115 3065
rect 5167 3013 5291 3065
rect 5343 3013 5467 3065
rect 5519 3013 6094 3065
rect 4577 3005 6094 3013
rect 5603 2711 6094 3005
rect 5603 2659 5630 2711
rect 5682 2659 5694 2711
rect 5746 2659 5758 2711
rect 5810 2659 5822 2711
rect 5874 2659 5886 2711
rect 5938 2659 5950 2711
rect 6002 2659 6014 2711
rect 6066 2659 6094 2711
rect -646 -603 -96 -486
rect -646 -2511 -452 -603
rect -208 -2511 -96 -603
rect 5603 -1754 6094 2659
rect 5603 -1806 5631 -1754
rect 5683 -1806 5695 -1754
rect 5747 -1806 5759 -1754
rect 5811 -1806 5823 -1754
rect 5875 -1806 5887 -1754
rect 5939 -1806 5951 -1754
rect 6003 -1806 6015 -1754
rect 6067 -1806 6094 -1754
rect 5603 -1814 6094 -1806
rect -646 -2615 -96 -2511
<< via2 >>
rect -49 3731 407 3947
rect -438 -2505 -222 -609
<< metal3 >>
rect -478 3951 594 4003
rect -478 3727 -53 3951
rect 411 3727 594 3951
rect -478 3673 594 3727
rect -646 -605 -96 -486
rect -646 -2509 -442 -605
rect -218 -2509 -96 -605
rect -646 -2615 -96 -2509
<< via3 >>
rect -53 3947 411 3951
rect -53 3731 -49 3947
rect -49 3731 407 3947
rect 407 3731 411 3947
rect -53 3727 411 3731
rect -442 -609 -218 -605
rect -442 -2505 -438 -609
rect -438 -2505 -222 -609
rect -222 -2505 -218 -609
rect -442 -2509 -218 -2505
<< metal4 >>
rect -1445 3951 1065 4016
rect -1445 3727 -53 3951
rect 411 3727 1065 3951
rect -1445 3672 1065 3727
rect -465 -488 -98 -486
rect -521 -605 -96 -488
rect -521 -639 -442 -605
rect -218 -639 -96 -605
rect -521 -875 -448 -639
rect -212 -875 -96 -639
rect -521 -959 -442 -875
rect -218 -959 -96 -875
rect -521 -1195 -448 -959
rect -212 -1195 -96 -959
rect -521 -1279 -442 -1195
rect -218 -1279 -96 -1195
rect -521 -1515 -448 -1279
rect -212 -1515 -96 -1279
rect -521 -1599 -442 -1515
rect -218 -1599 -96 -1515
rect -521 -1835 -448 -1599
rect -212 -1835 -96 -1599
rect -521 -1919 -442 -1835
rect -218 -1919 -96 -1835
rect -521 -2155 -448 -1919
rect -212 -2155 -96 -1919
rect -521 -2239 -442 -2155
rect -218 -2239 -96 -2155
rect -521 -2475 -448 -2239
rect -212 -2475 -96 -2239
rect -521 -2509 -442 -2475
rect -218 -2509 -96 -2475
rect -521 -2615 -96 -2509
<< via4 >>
rect -448 -875 -442 -639
rect -442 -875 -218 -639
rect -218 -875 -212 -639
rect -448 -1195 -442 -959
rect -442 -1195 -218 -959
rect -218 -1195 -212 -959
rect -448 -1515 -442 -1279
rect -442 -1515 -218 -1279
rect -218 -1515 -212 -1279
rect -448 -1835 -442 -1599
rect -442 -1835 -218 -1599
rect -218 -1835 -212 -1599
rect -448 -2155 -442 -1919
rect -442 -2155 -218 -1919
rect -218 -2155 -212 -1919
rect -448 -2475 -442 -2239
rect -442 -2475 -218 -2239
rect -218 -2475 -212 -2239
<< metal5 >>
rect -1254 -639 -98 -488
rect -1254 -875 -448 -639
rect -212 -875 -98 -639
rect -1254 -959 -98 -875
rect -1254 -1195 -448 -959
rect -212 -1195 -98 -959
rect -1254 -1279 -98 -1195
rect -1254 -1515 -448 -1279
rect -212 -1515 -98 -1279
rect -1254 -1599 -98 -1515
rect -1254 -1835 -448 -1599
rect -212 -1835 -98 -1599
rect -1254 -1919 -98 -1835
rect -1254 -2155 -448 -1919
rect -212 -2155 -98 -1919
rect -1254 -2239 -98 -2155
rect -1254 -2475 -448 -2239
rect -212 -2475 -98 -2239
rect -1254 -2615 -98 -2475
use sky130_fd_pr__nfet_01v8_lvt_C43HKJ  sky130_fd_pr__nfet_01v8_lvt_C43HKJ_0
timestamp 1640969486
transform 0 1 3692 -1 0 -1146
box -201 -940 201 940
use sky130_fd_pr__nfet_01v8_lvt_H2P3K4  sky130_fd_pr__nfet_01v8_lvt_H2P3K4_0
timestamp 1640969486
transform 0 1 1680 -1 0 -1146
box -201 -1000 201 1000
use sky130_fd_pr__res_high_po_0p35_A4PB2C  sky130_fd_pr__res_high_po_0p35_A4PB2C_0
timestamp 1640969486
transform 0 1 1431 -1 0 -1779
box -191 -638 191 638
use sky130_fd_pr__res_high_po_0p35_PGG99R  sky130_fd_pr__res_high_po_0p35_PGG99R_0
timestamp 1640969486
transform 0 1 2134 -1 0 -2310
box -191 -1588 191 1588
use ForwardAmp  ForwardAmp_0
timestamp 1640969486
transform 1 0 0 0 1 0
box 0 66 5705 5234
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_0
timestamp 1640969486
transform 0 -1 -3746 1 0 621
box -3351 -3101 3373 3101
use sky130_fd_pr__diode_pd2nw_05v5_WW7YB9  sky130_fd_pr__diode_pd2nw_05v5_WW7YB9_0
timestamp 1640969486
transform 1 0 151 0 1 -1251
box -466 -466 466 466
<< labels >>
rlabel metal1 s 4671 -1142 4671 -1142 4 VBIAS1
port 1 nsew
rlabel metal1 s 3743 -2313 3743 -2313 4 VBIAS2
port 2 nsew
rlabel metal1 s 2236 5234 2236 5234 4 VDD
port 3 nsew
rlabel metal1 s 2230 3010 2230 3010 4 S1
port 4 nsew
rlabel metal1 s 0 633 0 633 4 G2
port 5 nsew
<< end >>
