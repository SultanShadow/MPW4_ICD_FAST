magic
tech sky130A
magscale 1 2
timestamp 1640969486
<< nwell >>
rect -144 -662 144 662
<< pmoslvt >>
rect -50 -600 50 600
<< pdiff >>
rect -108 561 -50 600
rect -108 527 -96 561
rect -62 527 -50 561
rect -108 493 -50 527
rect -108 459 -96 493
rect -62 459 -50 493
rect -108 425 -50 459
rect -108 391 -96 425
rect -62 391 -50 425
rect -108 357 -50 391
rect -108 323 -96 357
rect -62 323 -50 357
rect -108 289 -50 323
rect -108 255 -96 289
rect -62 255 -50 289
rect -108 221 -50 255
rect -108 187 -96 221
rect -62 187 -50 221
rect -108 153 -50 187
rect -108 119 -96 153
rect -62 119 -50 153
rect -108 85 -50 119
rect -108 51 -96 85
rect -62 51 -50 85
rect -108 17 -50 51
rect -108 -17 -96 17
rect -62 -17 -50 17
rect -108 -51 -50 -17
rect -108 -85 -96 -51
rect -62 -85 -50 -51
rect -108 -119 -50 -85
rect -108 -153 -96 -119
rect -62 -153 -50 -119
rect -108 -187 -50 -153
rect -108 -221 -96 -187
rect -62 -221 -50 -187
rect -108 -255 -50 -221
rect -108 -289 -96 -255
rect -62 -289 -50 -255
rect -108 -323 -50 -289
rect -108 -357 -96 -323
rect -62 -357 -50 -323
rect -108 -391 -50 -357
rect -108 -425 -96 -391
rect -62 -425 -50 -391
rect -108 -459 -50 -425
rect -108 -493 -96 -459
rect -62 -493 -50 -459
rect -108 -527 -50 -493
rect -108 -561 -96 -527
rect -62 -561 -50 -527
rect -108 -600 -50 -561
rect 50 561 108 600
rect 50 527 62 561
rect 96 527 108 561
rect 50 493 108 527
rect 50 459 62 493
rect 96 459 108 493
rect 50 425 108 459
rect 50 391 62 425
rect 96 391 108 425
rect 50 357 108 391
rect 50 323 62 357
rect 96 323 108 357
rect 50 289 108 323
rect 50 255 62 289
rect 96 255 108 289
rect 50 221 108 255
rect 50 187 62 221
rect 96 187 108 221
rect 50 153 108 187
rect 50 119 62 153
rect 96 119 108 153
rect 50 85 108 119
rect 50 51 62 85
rect 96 51 108 85
rect 50 17 108 51
rect 50 -17 62 17
rect 96 -17 108 17
rect 50 -51 108 -17
rect 50 -85 62 -51
rect 96 -85 108 -51
rect 50 -119 108 -85
rect 50 -153 62 -119
rect 96 -153 108 -119
rect 50 -187 108 -153
rect 50 -221 62 -187
rect 96 -221 108 -187
rect 50 -255 108 -221
rect 50 -289 62 -255
rect 96 -289 108 -255
rect 50 -323 108 -289
rect 50 -357 62 -323
rect 96 -357 108 -323
rect 50 -391 108 -357
rect 50 -425 62 -391
rect 96 -425 108 -391
rect 50 -459 108 -425
rect 50 -493 62 -459
rect 96 -493 108 -459
rect 50 -527 108 -493
rect 50 -561 62 -527
rect 96 -561 108 -527
rect 50 -600 108 -561
<< pdiffc >>
rect -96 527 -62 561
rect -96 459 -62 493
rect -96 391 -62 425
rect -96 323 -62 357
rect -96 255 -62 289
rect -96 187 -62 221
rect -96 119 -62 153
rect -96 51 -62 85
rect -96 -17 -62 17
rect -96 -85 -62 -51
rect -96 -153 -62 -119
rect -96 -221 -62 -187
rect -96 -289 -62 -255
rect -96 -357 -62 -323
rect -96 -425 -62 -391
rect -96 -493 -62 -459
rect -96 -561 -62 -527
rect 62 527 96 561
rect 62 459 96 493
rect 62 391 96 425
rect 62 323 96 357
rect 62 255 96 289
rect 62 187 96 221
rect 62 119 96 153
rect 62 51 96 85
rect 62 -17 96 17
rect 62 -85 96 -51
rect 62 -153 96 -119
rect 62 -221 96 -187
rect 62 -289 96 -255
rect 62 -357 96 -323
rect 62 -425 96 -391
rect 62 -493 96 -459
rect 62 -561 96 -527
<< poly >>
rect -50 600 50 626
rect -50 -626 50 -600
<< locali >>
rect -96 561 -62 604
rect -96 493 -62 523
rect -96 425 -62 451
rect -96 357 -62 379
rect -96 289 -62 307
rect -96 221 -62 235
rect -96 153 -62 163
rect -96 85 -62 91
rect -96 17 -62 19
rect -96 -19 -62 -17
rect -96 -91 -62 -85
rect -96 -163 -62 -153
rect -96 -235 -62 -221
rect -96 -307 -62 -289
rect -96 -379 -62 -357
rect -96 -451 -62 -425
rect -96 -523 -62 -493
rect -96 -604 -62 -561
rect 62 561 96 604
rect 62 493 96 523
rect 62 425 96 451
rect 62 357 96 379
rect 62 289 96 307
rect 62 221 96 235
rect 62 153 96 163
rect 62 85 96 91
rect 62 17 96 19
rect 62 -19 96 -17
rect 62 -91 96 -85
rect 62 -163 96 -153
rect 62 -235 96 -221
rect 62 -307 96 -289
rect 62 -379 96 -357
rect 62 -451 96 -425
rect 62 -523 96 -493
rect 62 -604 96 -561
<< viali >>
rect -96 527 -62 557
rect -96 523 -62 527
rect -96 459 -62 485
rect -96 451 -62 459
rect -96 391 -62 413
rect -96 379 -62 391
rect -96 323 -62 341
rect -96 307 -62 323
rect -96 255 -62 269
rect -96 235 -62 255
rect -96 187 -62 197
rect -96 163 -62 187
rect -96 119 -62 125
rect -96 91 -62 119
rect -96 51 -62 53
rect -96 19 -62 51
rect -96 -51 -62 -19
rect -96 -53 -62 -51
rect -96 -119 -62 -91
rect -96 -125 -62 -119
rect -96 -187 -62 -163
rect -96 -197 -62 -187
rect -96 -255 -62 -235
rect -96 -269 -62 -255
rect -96 -323 -62 -307
rect -96 -341 -62 -323
rect -96 -391 -62 -379
rect -96 -413 -62 -391
rect -96 -459 -62 -451
rect -96 -485 -62 -459
rect -96 -527 -62 -523
rect -96 -557 -62 -527
rect 62 527 96 557
rect 62 523 96 527
rect 62 459 96 485
rect 62 451 96 459
rect 62 391 96 413
rect 62 379 96 391
rect 62 323 96 341
rect 62 307 96 323
rect 62 255 96 269
rect 62 235 96 255
rect 62 187 96 197
rect 62 163 96 187
rect 62 119 96 125
rect 62 91 96 119
rect 62 51 96 53
rect 62 19 96 51
rect 62 -51 96 -19
rect 62 -53 96 -51
rect 62 -119 96 -91
rect 62 -125 96 -119
rect 62 -187 96 -163
rect 62 -197 96 -187
rect 62 -255 96 -235
rect 62 -269 96 -255
rect 62 -323 96 -307
rect 62 -341 96 -323
rect 62 -391 96 -379
rect 62 -413 96 -391
rect 62 -459 96 -451
rect 62 -485 96 -459
rect 62 -527 96 -523
rect 62 -557 96 -527
<< metal1 >>
rect -102 557 -56 600
rect -102 523 -96 557
rect -62 523 -56 557
rect -102 485 -56 523
rect -102 451 -96 485
rect -62 451 -56 485
rect -102 413 -56 451
rect -102 379 -96 413
rect -62 379 -56 413
rect -102 341 -56 379
rect -102 307 -96 341
rect -62 307 -56 341
rect -102 269 -56 307
rect -102 235 -96 269
rect -62 235 -56 269
rect -102 197 -56 235
rect -102 163 -96 197
rect -62 163 -56 197
rect -102 125 -56 163
rect -102 91 -96 125
rect -62 91 -56 125
rect -102 53 -56 91
rect -102 19 -96 53
rect -62 19 -56 53
rect -102 -19 -56 19
rect -102 -53 -96 -19
rect -62 -53 -56 -19
rect -102 -91 -56 -53
rect -102 -125 -96 -91
rect -62 -125 -56 -91
rect -102 -163 -56 -125
rect -102 -197 -96 -163
rect -62 -197 -56 -163
rect -102 -235 -56 -197
rect -102 -269 -96 -235
rect -62 -269 -56 -235
rect -102 -307 -56 -269
rect -102 -341 -96 -307
rect -62 -341 -56 -307
rect -102 -379 -56 -341
rect -102 -413 -96 -379
rect -62 -413 -56 -379
rect -102 -451 -56 -413
rect -102 -485 -96 -451
rect -62 -485 -56 -451
rect -102 -523 -56 -485
rect -102 -557 -96 -523
rect -62 -557 -56 -523
rect -102 -600 -56 -557
rect 56 557 102 600
rect 56 523 62 557
rect 96 523 102 557
rect 56 485 102 523
rect 56 451 62 485
rect 96 451 102 485
rect 56 413 102 451
rect 56 379 62 413
rect 96 379 102 413
rect 56 341 102 379
rect 56 307 62 341
rect 96 307 102 341
rect 56 269 102 307
rect 56 235 62 269
rect 96 235 102 269
rect 56 197 102 235
rect 56 163 62 197
rect 96 163 102 197
rect 56 125 102 163
rect 56 91 62 125
rect 96 91 102 125
rect 56 53 102 91
rect 56 19 62 53
rect 96 19 102 53
rect 56 -19 102 19
rect 56 -53 62 -19
rect 96 -53 102 -19
rect 56 -91 102 -53
rect 56 -125 62 -91
rect 96 -125 102 -91
rect 56 -163 102 -125
rect 56 -197 62 -163
rect 96 -197 102 -163
rect 56 -235 102 -197
rect 56 -269 62 -235
rect 96 -269 102 -235
rect 56 -307 102 -269
rect 56 -341 62 -307
rect 96 -341 102 -307
rect 56 -379 102 -341
rect 56 -413 62 -379
rect 96 -413 102 -379
rect 56 -451 102 -413
rect 56 -485 62 -451
rect 96 -485 102 -451
rect 56 -523 102 -485
rect 56 -557 62 -523
rect 96 -557 102 -523
rect 56 -600 102 -557
<< end >>
