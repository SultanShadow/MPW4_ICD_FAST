magic
tech sky130A
magscale 1 2
timestamp 1640969486
<< nwell >>
rect 1289 562 2686 564
rect -917 558 2686 562
rect -1693 549 2686 558
rect -3322 -373 2686 549
rect -3322 -377 1315 -373
rect -3322 -379 4 -377
rect -3322 -380 -3120 -379
<< poly >>
rect -2894 462 2337 482
rect -2894 428 -2844 462
rect -2810 428 -2776 462
rect -2742 428 -2708 462
rect -2674 428 -2640 462
rect -2606 428 -2572 462
rect -2538 428 -2504 462
rect -2470 428 -2436 462
rect -2402 428 -2368 462
rect -2334 428 -2300 462
rect -2266 428 -2232 462
rect -2198 428 -2164 462
rect -2130 428 -2096 462
rect -2062 428 -2028 462
rect -1994 428 -1960 462
rect -1926 428 -1892 462
rect -1858 428 -1824 462
rect -1790 428 -1756 462
rect -1722 428 -1688 462
rect -1654 428 -1620 462
rect -1586 428 -1552 462
rect -1518 428 -1484 462
rect -1450 428 -1416 462
rect -1382 428 -1348 462
rect -1314 428 -1280 462
rect -1246 428 -1212 462
rect -1178 428 -1144 462
rect -1110 428 -1076 462
rect -1042 428 -1008 462
rect -974 428 -940 462
rect -906 428 -872 462
rect -838 428 -804 462
rect -770 428 -736 462
rect -702 428 -668 462
rect -634 428 -600 462
rect -566 428 -532 462
rect -498 428 -464 462
rect -430 428 -396 462
rect -362 428 -328 462
rect -294 428 -260 462
rect -226 428 -192 462
rect -158 428 -124 462
rect -90 428 -56 462
rect -22 428 12 462
rect 46 428 80 462
rect 114 428 148 462
rect 182 428 216 462
rect 250 428 284 462
rect 318 428 352 462
rect 386 428 420 462
rect 454 428 488 462
rect 522 428 556 462
rect 590 428 624 462
rect 658 428 692 462
rect 726 428 760 462
rect 794 428 828 462
rect 862 428 896 462
rect 930 428 964 462
rect 998 428 1032 462
rect 1066 428 1100 462
rect 1134 428 1168 462
rect 1202 428 1236 462
rect 1270 428 1304 462
rect 1338 428 1372 462
rect 1406 428 1440 462
rect 1474 428 1508 462
rect 1542 428 1576 462
rect 1610 428 1644 462
rect 1678 428 1712 462
rect 1746 428 1780 462
rect 1814 428 1848 462
rect 1882 428 1916 462
rect 1950 428 1984 462
rect 2018 428 2052 462
rect 2086 428 2120 462
rect 2154 428 2188 462
rect 2222 428 2256 462
rect 2290 428 2337 462
rect -2894 407 2337 428
rect -2894 404 2338 407
rect -2894 311 -1894 404
rect -1836 311 -836 404
rect -778 311 222 404
rect 280 311 1280 404
rect 1338 311 2338 404
<< polycont >>
rect -2844 428 -2810 462
rect -2776 428 -2742 462
rect -2708 428 -2674 462
rect -2640 428 -2606 462
rect -2572 428 -2538 462
rect -2504 428 -2470 462
rect -2436 428 -2402 462
rect -2368 428 -2334 462
rect -2300 428 -2266 462
rect -2232 428 -2198 462
rect -2164 428 -2130 462
rect -2096 428 -2062 462
rect -2028 428 -1994 462
rect -1960 428 -1926 462
rect -1892 428 -1858 462
rect -1824 428 -1790 462
rect -1756 428 -1722 462
rect -1688 428 -1654 462
rect -1620 428 -1586 462
rect -1552 428 -1518 462
rect -1484 428 -1450 462
rect -1416 428 -1382 462
rect -1348 428 -1314 462
rect -1280 428 -1246 462
rect -1212 428 -1178 462
rect -1144 428 -1110 462
rect -1076 428 -1042 462
rect -1008 428 -974 462
rect -940 428 -906 462
rect -872 428 -838 462
rect -804 428 -770 462
rect -736 428 -702 462
rect -668 428 -634 462
rect -600 428 -566 462
rect -532 428 -498 462
rect -464 428 -430 462
rect -396 428 -362 462
rect -328 428 -294 462
rect -260 428 -226 462
rect -192 428 -158 462
rect -124 428 -90 462
rect -56 428 -22 462
rect 12 428 46 462
rect 80 428 114 462
rect 148 428 182 462
rect 216 428 250 462
rect 284 428 318 462
rect 352 428 386 462
rect 420 428 454 462
rect 488 428 522 462
rect 556 428 590 462
rect 624 428 658 462
rect 692 428 726 462
rect 760 428 794 462
rect 828 428 862 462
rect 896 428 930 462
rect 964 428 998 462
rect 1032 428 1066 462
rect 1100 428 1134 462
rect 1168 428 1202 462
rect 1236 428 1270 462
rect 1304 428 1338 462
rect 1372 428 1406 462
rect 1440 428 1474 462
rect 1508 428 1542 462
rect 1576 428 1610 462
rect 1644 428 1678 462
rect 1712 428 1746 462
rect 1780 428 1814 462
rect 1848 428 1882 462
rect 1916 428 1950 462
rect 1984 428 2018 462
rect 2052 428 2086 462
rect 2120 428 2154 462
rect 2188 428 2222 462
rect 2256 428 2290 462
<< locali >>
rect -2894 462 2337 482
rect -2894 428 -2851 462
rect -2810 428 -2779 462
rect -2742 428 -2708 462
rect -2673 428 -2640 462
rect -2601 428 -2572 462
rect -2529 428 -2504 462
rect -2457 428 -2436 462
rect -2385 428 -2368 462
rect -2313 428 -2300 462
rect -2241 428 -2232 462
rect -2169 428 -2164 462
rect -2097 428 -2096 462
rect -2062 428 -2059 462
rect -1994 428 -1987 462
rect -1926 428 -1915 462
rect -1858 428 -1843 462
rect -1790 428 -1771 462
rect -1722 428 -1699 462
rect -1654 428 -1627 462
rect -1586 428 -1555 462
rect -1518 428 -1484 462
rect -1449 428 -1416 462
rect -1377 428 -1348 462
rect -1305 428 -1280 462
rect -1233 428 -1212 462
rect -1161 428 -1144 462
rect -1089 428 -1076 462
rect -1017 428 -1008 462
rect -945 428 -940 462
rect -873 428 -872 462
rect -838 428 -835 462
rect -770 428 -763 462
rect -702 428 -691 462
rect -634 428 -619 462
rect -566 428 -547 462
rect -498 428 -475 462
rect -430 428 -403 462
rect -362 428 -331 462
rect -294 428 -260 462
rect -225 428 -192 462
rect -153 428 -124 462
rect -81 428 -56 462
rect -9 428 12 462
rect 63 428 80 462
rect 135 428 148 462
rect 207 428 216 462
rect 279 428 284 462
rect 351 428 352 462
rect 386 428 389 462
rect 454 428 461 462
rect 522 428 533 462
rect 590 428 605 462
rect 658 428 677 462
rect 726 428 749 462
rect 794 428 821 462
rect 862 428 893 462
rect 930 428 964 462
rect 999 428 1032 462
rect 1071 428 1100 462
rect 1143 428 1168 462
rect 1215 428 1236 462
rect 1287 428 1304 462
rect 1359 428 1372 462
rect 1431 428 1440 462
rect 1503 428 1508 462
rect 1575 428 1576 462
rect 1610 428 1613 462
rect 1678 428 1685 462
rect 1746 428 1757 462
rect 1814 428 1829 462
rect 1882 428 1901 462
rect 1950 428 1973 462
rect 2018 428 2045 462
rect 2086 428 2117 462
rect 2154 428 2188 462
rect 2223 428 2256 462
rect 2295 428 2337 462
rect -2894 402 2337 428
rect -2939 -173 -2905 -118
rect -823 -173 -789 -118
rect 1293 -173 1327 -118
rect -2939 -217 1328 -173
<< viali >>
rect -2851 428 -2844 462
rect -2844 428 -2817 462
rect -2779 428 -2776 462
rect -2776 428 -2745 462
rect -2707 428 -2674 462
rect -2674 428 -2673 462
rect -2635 428 -2606 462
rect -2606 428 -2601 462
rect -2563 428 -2538 462
rect -2538 428 -2529 462
rect -2491 428 -2470 462
rect -2470 428 -2457 462
rect -2419 428 -2402 462
rect -2402 428 -2385 462
rect -2347 428 -2334 462
rect -2334 428 -2313 462
rect -2275 428 -2266 462
rect -2266 428 -2241 462
rect -2203 428 -2198 462
rect -2198 428 -2169 462
rect -2131 428 -2130 462
rect -2130 428 -2097 462
rect -2059 428 -2028 462
rect -2028 428 -2025 462
rect -1987 428 -1960 462
rect -1960 428 -1953 462
rect -1915 428 -1892 462
rect -1892 428 -1881 462
rect -1843 428 -1824 462
rect -1824 428 -1809 462
rect -1771 428 -1756 462
rect -1756 428 -1737 462
rect -1699 428 -1688 462
rect -1688 428 -1665 462
rect -1627 428 -1620 462
rect -1620 428 -1593 462
rect -1555 428 -1552 462
rect -1552 428 -1521 462
rect -1483 428 -1450 462
rect -1450 428 -1449 462
rect -1411 428 -1382 462
rect -1382 428 -1377 462
rect -1339 428 -1314 462
rect -1314 428 -1305 462
rect -1267 428 -1246 462
rect -1246 428 -1233 462
rect -1195 428 -1178 462
rect -1178 428 -1161 462
rect -1123 428 -1110 462
rect -1110 428 -1089 462
rect -1051 428 -1042 462
rect -1042 428 -1017 462
rect -979 428 -974 462
rect -974 428 -945 462
rect -907 428 -906 462
rect -906 428 -873 462
rect -835 428 -804 462
rect -804 428 -801 462
rect -763 428 -736 462
rect -736 428 -729 462
rect -691 428 -668 462
rect -668 428 -657 462
rect -619 428 -600 462
rect -600 428 -585 462
rect -547 428 -532 462
rect -532 428 -513 462
rect -475 428 -464 462
rect -464 428 -441 462
rect -403 428 -396 462
rect -396 428 -369 462
rect -331 428 -328 462
rect -328 428 -297 462
rect -259 428 -226 462
rect -226 428 -225 462
rect -187 428 -158 462
rect -158 428 -153 462
rect -115 428 -90 462
rect -90 428 -81 462
rect -43 428 -22 462
rect -22 428 -9 462
rect 29 428 46 462
rect 46 428 63 462
rect 101 428 114 462
rect 114 428 135 462
rect 173 428 182 462
rect 182 428 207 462
rect 245 428 250 462
rect 250 428 279 462
rect 317 428 318 462
rect 318 428 351 462
rect 389 428 420 462
rect 420 428 423 462
rect 461 428 488 462
rect 488 428 495 462
rect 533 428 556 462
rect 556 428 567 462
rect 605 428 624 462
rect 624 428 639 462
rect 677 428 692 462
rect 692 428 711 462
rect 749 428 760 462
rect 760 428 783 462
rect 821 428 828 462
rect 828 428 855 462
rect 893 428 896 462
rect 896 428 927 462
rect 965 428 998 462
rect 998 428 999 462
rect 1037 428 1066 462
rect 1066 428 1071 462
rect 1109 428 1134 462
rect 1134 428 1143 462
rect 1181 428 1202 462
rect 1202 428 1215 462
rect 1253 428 1270 462
rect 1270 428 1287 462
rect 1325 428 1338 462
rect 1338 428 1359 462
rect 1397 428 1406 462
rect 1406 428 1431 462
rect 1469 428 1474 462
rect 1474 428 1503 462
rect 1541 428 1542 462
rect 1542 428 1575 462
rect 1613 428 1644 462
rect 1644 428 1647 462
rect 1685 428 1712 462
rect 1712 428 1719 462
rect 1757 428 1780 462
rect 1780 428 1791 462
rect 1829 428 1848 462
rect 1848 428 1863 462
rect 1901 428 1916 462
rect 1916 428 1935 462
rect 1973 428 1984 462
rect 1984 428 2007 462
rect 2045 428 2052 462
rect 2052 428 2079 462
rect 2117 428 2120 462
rect 2120 428 2151 462
rect 2189 428 2222 462
rect 2222 428 2223 462
rect 2261 428 2290 462
rect 2290 428 2295 462
<< metal1 >>
rect -2894 462 2337 482
rect -2894 428 -2851 462
rect -2817 428 -2779 462
rect -2745 428 -2707 462
rect -2673 428 -2635 462
rect -2601 428 -2563 462
rect -2529 428 -2491 462
rect -2457 428 -2419 462
rect -2385 428 -2347 462
rect -2313 428 -2275 462
rect -2241 428 -2203 462
rect -2169 428 -2131 462
rect -2097 428 -2059 462
rect -2025 428 -1987 462
rect -1953 428 -1915 462
rect -1881 428 -1843 462
rect -1809 428 -1771 462
rect -1737 428 -1699 462
rect -1665 428 -1627 462
rect -1593 428 -1555 462
rect -1521 428 -1483 462
rect -1449 428 -1411 462
rect -1377 428 -1339 462
rect -1305 428 -1267 462
rect -1233 428 -1195 462
rect -1161 428 -1123 462
rect -1089 428 -1051 462
rect -1017 428 -979 462
rect -945 428 -907 462
rect -873 428 -835 462
rect -801 428 -763 462
rect -729 428 -691 462
rect -657 428 -619 462
rect -585 428 -547 462
rect -513 428 -475 462
rect -441 428 -403 462
rect -369 428 -331 462
rect -297 428 -259 462
rect -225 428 -187 462
rect -153 428 -115 462
rect -81 428 -43 462
rect -9 428 29 462
rect 63 428 101 462
rect 135 428 173 462
rect 207 428 245 462
rect 279 428 317 462
rect 351 428 389 462
rect 423 428 461 462
rect 495 428 533 462
rect 567 428 605 462
rect 639 428 677 462
rect 711 428 749 462
rect 783 428 821 462
rect 855 428 893 462
rect 927 428 965 462
rect 999 428 1037 462
rect 1071 428 1109 462
rect 1143 428 1181 462
rect 1215 428 1253 462
rect 1287 428 1325 462
rect 1359 428 1397 462
rect 1431 428 1469 462
rect 1503 428 1541 462
rect 1575 428 1613 462
rect 1647 428 1685 462
rect 1719 428 1757 462
rect 1791 428 1829 462
rect 1863 428 1901 462
rect 1935 428 1973 462
rect 2007 428 2045 462
rect 2079 428 2117 462
rect 2151 428 2189 462
rect 2223 428 2261 462
rect 2295 428 2337 462
rect -2894 402 2337 428
rect -1881 -181 -1847 -97
rect 235 -143 269 -97
rect 234 -181 269 -143
rect 2351 -181 2385 -97
rect -1882 -184 2385 -181
rect -1882 -218 2384 -184
use sky130_fd_pr__pfet_g5v0d10v5_9HRSSM  sky130_fd_pr__pfet_g5v0d10v5_9HRSSM_4
timestamp 1640969486
transform 1 0 1839 0 1 85
box -624 -266 624 266
use sky130_fd_pr__pfet_g5v0d10v5_9HRSSM  sky130_fd_pr__pfet_g5v0d10v5_9HRSSM_3
timestamp 1640969486
transform 1 0 781 0 1 85
box -624 -266 624 266
use sky130_fd_pr__pfet_g5v0d10v5_9HRSSM  sky130_fd_pr__pfet_g5v0d10v5_9HRSSM_2
timestamp 1640969486
transform 1 0 -277 0 1 85
box -624 -266 624 266
use sky130_fd_pr__pfet_g5v0d10v5_9HRSSM  sky130_fd_pr__pfet_g5v0d10v5_9HRSSM_1
timestamp 1640969486
transform 1 0 -1335 0 1 85
box -624 -266 624 266
use sky130_fd_pr__pfet_g5v0d10v5_9HRSSM  sky130_fd_pr__pfet_g5v0d10v5_9HRSSM_0
timestamp 1640969486
transform 1 0 -2393 0 1 85
box -624 -266 624 266
<< labels >>
flabel locali s -2619 -207 -2619 -207 0 FreeSans 2500 0 0 0 S
port 1 nsew
flabel metal1 s 1786 -207 1786 -207 0 FreeSans 2500 0 0 0 D
port 2 nsew
flabel locali s 35 434 35 434 0 FreeSans 2500 0 0 0 G
port 3 nsew
<< end >>
